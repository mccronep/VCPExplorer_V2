netcdf raob_oun-20040520_1200 {
dimensions:
	recNum = UNLIMITED ; // (134 currently)
	manLevel = 22 ;
	sigTLevel = 150 ;
	sigWLevel = 76 ;
	mWndNum = 4 ;
	mTropNum = 4 ;
	staNameLen = 50 ;
	maxStaticIds = 500 ;
	totalIdLen = 50 ;
	nInventoryBins = 32 ;
variables:
	int nStaticIds ;
		nStaticIds:_FillValue = 0 ;
	char staticIds(maxStaticIds, totalIdLen) ;
		staticIds:_FillValue = "" ;
	int lastRecord(maxStaticIds) ;
		lastRecord:_FillValue = -1 ;
	int invTime(recNum) ;
		invTime:_FillValue = 0 ;
	int prevRecord(recNum) ;
		prevRecord:_FillValue = -1 ;
	int inventory(maxStaticIds) ;
		inventory:_FillValue = 0 ;
	int globalInventory ;
		globalInventory:_FillValue = 0 ;
	int firstOverflow ;
		firstOverflow:_FillValue = -1 ;
	int isOverflow(recNum) ;
		isOverflow:_FillValue = 0 ;
	int firstInBin(nInventoryBins) ;
		firstInBin:_FillValue = -1 ;
	int lastInBin(nInventoryBins) ;
		lastInBin:_FillValue = -1 ;
	int wmoStaNum(recNum) ;
		wmoStaNum:long_name = "WMO Station Number" ;
		wmoStaNum:reference = "Volume A of WMO publication 9" ;
		wmoStaNum:_FillValue = 99999 ;
	char staName(recNum, staNameLen) ;
		staName:long_name = "Station Identifier" ;
	float staLat(recNum) ;
		staLat:long_name = "Station Latitude" ;
		staLat:units = "degree_N" ;
		staLat:valid_range = 0.f, 90.f ;
		staLat:_FillValue = 99999.f ;
	float staLon(recNum) ;
		staLon:long_name = "Station Longitude" ;
		staLon:units = "degree_E" ;
		staLon:valid_range = -180.f, -50.f ;
		staLon:_FillValue = 99999.f ;
	float staElev(recNum) ;
		staElev:long_name = "Station Elevation" ;
		staElev:units = "meter" ;
		staElev:valid_range = -100.f, 3500.f ;
		staElev:_FillValue = 99999.f ;
	double synTime(recNum) ;
		synTime:long_name = "Synoptic Time" ;
		synTime:units = "seconds since (1970-1-1 00:00:0.0)" ;
	int numMand(recNum) ;
		numMand:long_name = "Number of Mandatory Levels" ;
		numMand:valid_range = 0, 22 ;
		numMand:_FillValue = 99999 ;
	int numSigT(recNum) ;
		numSigT:long_name = "Number of Significant Levels wrt T" ;
		numSigT:valid_range = 0, 150 ;
		numSigT:_FillValue = 99999 ;
	int numSigW(recNum) ;
		numSigW:long_name = "Number of Significant Levels wrt W" ;
		numSigW:valid_range = 0, 76 ;
		numSigW:_FillValue = 99999 ;
	int numMwnd(recNum) ;
		numMwnd:long_name = "Number of Maximum Wind Levels" ;
		numMwnd:valid_range = 0, 4 ;
		numMwnd:_FillValue = 99999 ;
	int numTrop(recNum) ;
		numTrop:long_name = "Number of Tropopause Levels" ;
		numTrop:valid_range = 0, 4 ;
		numTrop:_FillValue = 99999 ;
	double relTime(recNum) ;
		relTime:long_name = "Sounding Release Time" ;
		relTime:units = "seconds since (1970-1-1 00:00:0.0)" ;
		relTime:_FillValue = -1.e+38 ;
	int sondTyp(recNum) ;
		sondTyp:long_name = "Instrument Type" ;
		sondTyp:reference = "Federal Meteorological Handbook No. 4" ;
		sondTyp:_FillValue = 99999 ;
	float prMan(recNum, manLevel) ;
		prMan:long_name = "Pressure - Mandatory level" ;
		prMan:units = "hectopascal" ;
		prMan:valid_range = 1.f, 1500.f ;
		prMan:_FillValue = 99999.f ;
	float htMan(recNum, manLevel) ;
		htMan:long_name = "Geopotential - Mandatory level" ;
		htMan:units = "meter" ;
		htMan:valid_range = -250.f, 60000.f ;
		htMan:_FillValue = 99999.f ;
	float tpMan(recNum, manLevel) ;
		tpMan:long_name = "Temperature - Mandatory level" ;
		tpMan:units = "kelvin" ;
		tpMan:valid_range = 173.f, 373.f ;
		tpMan:_FillValue = 99999.f ;
	float tdMan(recNum, manLevel) ;
		tdMan:long_name = "Dew Point Depression - Mandatory level" ;
		tdMan:units = "kelvin" ;
		tdMan:valid_range = 0.f, 60.f ;
		tdMan:_FillValue = 99999.f ;
	float wdMan(recNum, manLevel) ;
		wdMan:long_name = "Wind Direction - Mandatory level" ;
		wdMan:units = "degree_true" ;
		wdMan:valid_range = 0.f, 360.f ;
		wdMan:_FillValue = 99999.f ;
	float wsMan(recNum, manLevel) ;
		wsMan:long_name = "Wind Speed - Mandatory level" ;
		wsMan:units = "meter/sec" ;
		wsMan:valid_range = 0.f, 300.f ;
		wsMan:_FillValue = 99999.f ;
	float prSigT(recNum, sigTLevel) ;
		prSigT:long_name = "Pressure - Significant level wrt T" ;
		prSigT:units = "hectopascal" ;
		prSigT:valid_range = 1.f, 1500.f ;
		prSigT:_FillValue = 99999.f ;
	float tpSigT(recNum, sigTLevel) ;
		tpSigT:long_name = "Temperature - Significant level wrt T" ;
		tpSigT:units = "kelvin" ;
		tpSigT:valid_range = 173.f, 373.f ;
		tpSigT:_FillValue = 99999.f ;
	float tdSigT(recNum, sigTLevel) ;
		tdSigT:long_name = "Dew Point Depression - Significant level wrt T" ;
		tdSigT:units = "kelvin" ;
		tdSigT:valid_range = 0.f, 60.f ;
		tdSigT:_FillValue = 99999.f ;
	float htSigW(recNum, sigWLevel) ;
		htSigW:long_name = "Geopotential - Significant level wrt W" ;
		htSigW:units = "meter" ;
		htSigW:valid_range = -250.f, 60000.f ;
		htSigW:_FillValue = 99999.f ;
	float wdSigW(recNum, sigWLevel) ;
		wdSigW:long_name = "Wind Direction - Significant level wrt W" ;
		wdSigW:units = "degree_true" ;
		wdSigW:valid_range = 0.f, 360.f ;
		wdSigW:_FillValue = 99999.f ;
	float wsSigW(recNum, sigWLevel) ;
		wsSigW:long_name = "Wind Speed - Significant level wrt W" ;
		wsSigW:units = "meter/sec" ;
		wsSigW:valid_range = 0.f, 300.f ;
		wsSigW:_FillValue = 99999.f ;
	float prTrop(recNum, mTropNum) ;
		prTrop:long_name = "Pressure - Tropopause level" ;
		prTrop:units = "hectopascal" ;
		prTrop:valid_range = 1.f, 1500.f ;
		prTrop:_FillValue = 99999.f ;
	float tpTrop(recNum, mTropNum) ;
		tpTrop:long_name = "Temperature - Tropopause level" ;
		tpTrop:units = "kelvin" ;
		tpTrop:valid_range = 173.f, 373.f ;
		tpTrop:_FillValue = 99999.f ;
	float tdTrop(recNum, mTropNum) ;
		tdTrop:long_name = "Dew Point Depression - Tropopause level" ;
		tdTrop:units = "kelvin" ;
		tdTrop:valid_range = 0.f, 60.f ;
		tdTrop:_FillValue = 99999.f ;
	float wdTrop(recNum, mTropNum) ;
		wdTrop:long_name = "Wind Direction - Tropopause level" ;
		wdTrop:units = "degree_true" ;
		wdTrop:valid_range = 0.f, 360.f ;
		wdTrop:_FillValue = 99999.f ;
	float wsTrop(recNum, mTropNum) ;
		wsTrop:long_name = "Wind Speed - Tropopause level" ;
		wsTrop:units = "meter/sec" ;
		wsTrop:valid_range = 0.f, 300.f ;
		wsTrop:_FillValue = 99999.f ;
	float prMaxW(recNum, mWndNum) ;
		prMaxW:long_name = "Pressure - Maximum wind level" ;
		prMaxW:units = "hectopascal" ;
		prMaxW:valid_range = 1.f, 1500.f ;
		prMaxW:_FillValue = 99999.f ;
	float wdMaxW(recNum, mWndNum) ;
		wdMaxW:long_name = "Wind Direction - Maximum wind level" ;
		wdMaxW:units = "degree_true" ;
		wdMaxW:valid_range = 0.f, 360.f ;
		wdMaxW:_FillValue = 99999.f ;
	float wsMaxW(recNum, mWndNum) ;
		wsMaxW:long_name = "Wind Speed - Maximum wind level" ;
		wsMaxW:units = "meter/sec" ;
		wsMaxW:valid_range = 0.f, 300.f ;
		wsMaxW:_FillValue = 99999.f ;

// global attributes:
		:comment0 = "First mandatory level is surface level" ;
		:version = "Forecast Systems Lab 5.0" ;
		:cdlDate = "20000118" ;
		:idVariables = "staName" ;
		:timeVariables = "synTime" ;
		:latLonVars = "staLat,staLon" ;
		:filePeriod = 43200 ;
		:fileEndOffset = 43199 ;
data:

 nStaticIds = 133 ;

 staticIds =
  "7460",
  "CWEG",
  "CWEU",
  "CWMW",
  "CWPL",
  "CWSA",
  "CWZC",
  "CYBK",
  "CYCB",
  "CYEV",
  "CYFB",
  "CYJT",
  "CYLT",
  "CYLW",
  "CYPH",
  "CYQD",
  "CYQI",
  "CYRB",
  "CYSM",
  "CYUX",
  "CYVP",
  "CYVQ",
  "CYXY",
  "CYYE",
  "CYYR",
  "CYYT",
  "CYZT",
  "CYZV",
  "K1Y7",
  "KABQ",
  "KABR",
  "KALB",
  "KAMA",
  "KAPX",
  "KBIS",
  "KBMX",
  "KBOI",
  "KBRO",
  "KBUF",
  "KCAR",
  "KCHH",
  "KCHS",
  "KCRP",
  "KDDC",
  "KDNR",
  "KDRA",
  "KDRT",
  "KDTX",
  "KDVN",
  "KEDW",
  "KEPZ",
  "KEYW",
  "KFFC",
  "KFGZ",
  "KFWD",
  "KGGW",
  "KGJT",
  "KGRB",
  "KGSO",
  "KGYX",
  "KILN",
  "KILX",
  "KINL",
  "KJAN",
  "KJAX",
  "KLBF",
  "KLCH",
  "KLIX",
  "KLKN",
  "KLWX",
  "KLZK",
  "KMAF",
  "KMFL",
  "KMFR",
  "KMHX",
  "KMPX",
  "KNKX",
  "KNSI",
  "KOAK",
  "KOAX",
  "KOHX",
  "KOKX",
  "KOTX",
  "KOUN",
  "KPIT",
  "KREV",
  "KRIW",
  "KRNK",
  "KSGF",
  "KSHV",
  "KSLC",
  "KTBW",
  "KTFX",
  "KTLH",
  "KTUS",
  "KUIL",
  "KUNR",
  "KVBG",
  "KWAL",
  "MACC",
  "MKJP",
  "MYNN",
  "MZBZ",
  "NSTU",
  "NTMN",
  "PABE",
  "PABR",
  "PACB",
  "PADQ",
  "PAFA",
  "PAFC",
  "PAKN",
  "PAMC",
  "PANT",
  "PAOM",
  "PAOT",
  "PASN",
  "PASY",
  "PAYA",
  "PGAC",
  "PGUM",
  "PHLI",
  "PHTO",
  "PJON",
  "PKWA",
  "PMKJ",
  "PTKK",
  "PTPN",
  "PTRO",
  "PTYA",
  "RJAM",
  "TJSJ",
  "TXKF",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 lastRecord = 5, 124, 120, 73, 108, 119, 116, 30, 121, 113, 110, 74, 105, 
    118, 76, 109, 72, 111, 112, 71, 75, 115, 114, 7, 107, 29, 123, 106, 126, 
    53, 65, 38, 51, 96, 27, 15, 66, 89, 87, 41, 43, 80, 90, 57, 58, 55, 47, 
    40, 101, 130, 52, 78, 82, 54, 46, 68, 59, 64, 34, 42, 37, 44, 67, 32, 79, 
    62, 83, 45, 63, 77, 49, 48, 31, 95, 33, 97, 92, 129, 60, 61, 35, 86, 69, 
    50, 39, 93, 26, 85, 56, 84, 94, 25, 99, 81, 91, 100, 98, 4, 36, 117, 127, 
    1, 125, 28, 133, 17, 2, 10, 12, 19, 20, 11, 18, 22, 8, 16, 9, 128, 21, 
    131, 70, 13, 23, 132, 104, 102, 24, 6, 14, 103, 122, 88, 0, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 invTime = 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085058000, 1085058000, 
    1085054400, 1085054400, 1085054400 ;

 prevRecord = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 3, _, _, _ ;

 inventory = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 5, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 globalInventory = 5 ;

 firstOverflow = _ ;

 isOverflow = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 firstInBin = 0, _, 129, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _ ;

 lastInBin = 133, _, 130, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _ ;

 wmoStaNum = 78016, 78073, 70026, 72381, 72393, 74606, 91348, 71945, 70200, 
    70308, 70316, 70326, 70350, 91165, 91408, 72230, 70133, 70219, 70231, 
    70261, 70273, 70361, 70398, 91285, 91334, 72210, 72672, 72764, 91765, 
    71801, 71926, 72202, 72235, 72305, 72317, 72327, 72402, 72426, 72518, 
    72520, 72632, 72712, 74389, 74494, 74560, 72233, 72249, 72261, 72265, 
    72340, 72357, 72363, 72364, 72365, 72376, 72387, 72440, 72451, 72469, 
    72476, 72493, 72558, 72562, 72582, 72645, 72659, 72681, 72747, 72768, 
    72786, 91212, 71081, 71603, 71722, 71815, 71906, 71907, 72403, 72201, 
    72206, 72208, 72214, 72215, 72240, 72248, 72318, 72501, 72528, 78526, 
    72250, 72251, 72274, 72293, 72489, 72572, 72597, 72634, 72649, 72662, 
    72776, 72797, 74455, 91376, 91413, 91366, 71082, 71811, 71816, 71845, 
    71867, 71909, 71924, 71934, 71957, 71964, 71043, 71836, 78988, 71203, 
    71600, 71917, 71925, 47991, 71109, 71119, 78583, 74004, 78397, 70414, 
    72291, 72381, 91217, 91275, 91925 ;

 staName =
  "TXKF",
  "MYNN",
  "PABR",
  "KEDW",
  "KVBG",
  "7460",
  "PTPN",
  "CYYE",
  "PAOM",
  "PASN",
  "PACB",
  "PAKN",
  "PADQ",
  "PHLI",
  "PTRO",
  "KBMX",
  "PAOT",
  "PABE",
  "PAMC",
  "PAFA",
  "PAFC",
  "PAYA",
  "PANT",
  "PHTO",
  "PTKK",
  "KTBW",
  "KRIW",
  "KBIS",
  "NSTU",
  "CYYT",
  "CYBK",
  "KMFL",
  "KJAN",
  "KMHX",
  "KGSO",
  "KOHX",
  "KWAL",
  "KILN",
  "KALB",
  "KPIT",
  "KDTX",
  "KCAR",
  "KGYX",
  "KCHH",
  "KILX",
  "KLIX",
  "KFWD",
  "KDRT",
  "KMAF",
  "KLZK",
  "KOUN",
  "KAMA",
  "KEPZ",
  "KABQ",
  "KFGZ",
  "KDRA",
  "KSGF",
  "KDDC",
  "KDNR",
  "KGJT",
  "KOAK",
  "KOAX",
  "KLBF",
  "KLKN",
  "KGRB",
  "KABR",
  "KBOI",
  "KINL",
  "KGGW",
  "KOTX",
  "PGUM",
  "CYUX",
  "CYQI",
  "CWMW",
  "CYJT",
  "CYVP",
  "CYPH",
  "KLWX",
  "KEYW",
  "KJAX",
  "KCHS",
  "KTLH",
  "KFFC",
  "KLCH",
  "KSHV",
  "KRNK",
  "KOKX",
  "KBUF",
  "TJSJ",
  "KBRO",
  "KCRP",
  "KTUS",
  "KNKX",
  "KREV",
  "KSLC",
  "KMFR",
  "KAPX",
  "KMPX",
  "KUNR",
  "KTFX",
  "KUIL",
  "KDVN",
  "PMKJ",
  "PTYA",
  "PKWA",
  "CYLT",
  "CYZV",
  "CYYR",
  "CWPL",
  "CYQD",
  "CYFB",
  "CYRB",
  "CYSM",
  "CYEV",
  "CYXY",
  "CYVQ",
  "CWZC",
  "MACC",
  "CYLW",
  "CWSA",
  "CWEU",
  "CYCB",
  "RJAM",
  "CYZT",
  "CWEG",
  "MZBZ",
  "K1Y7",
  "MKJP",
  "PASY",
  "KNSI",
  "KEDW",
  "PGAC",
  "PJON",
  "NTMN" ;

 staLat = 32.36667, 25.05, 71.28833, 34.93, 34.76, 34.65, 6.96667, 58.84, 
    64.51528, 57.11667, 55.20806, 58.67944, 57.75, 21.98333, 7.33333, 
    33.18028, 66.86667, 60.78333, 62.96667, 64.81528, 61.15694, 59.50801, 
    55.03944, 19.71667, 7.45528, 27.705, 43.06472, 46.77194, -14.33333, 
    47.68, 64.3, 25.75472, 32.32028, 34.77556, 36.08333, 36.23333, 37.93333, 
    39.42111, 42.73333, 40.53194, 42.69917, 46.86667, 43.8925, 41.66667, 
    40.15111, 30.33889, 32.835, 29.36667, 31.94278, 34.83556, 35.23556, 
    35.23194, 31.8775, 35.03806, 35.23056, 36.62861, 37.23583, 37.76139, 
    39.76806, 39.11667, 37.74306, 41.31944, 41.14972, 40.86028, 44.48889, 
    45.45444, 43.58, 48.56444, 48.20583, 47.68111, 13.47889, 68.78, 43.84, 
    46.39, 48.54, 58.11, 58.46, 38.98333, 24.55, 30.48472, 32.90056, 
    30.39583, 33.35583, 30.12528, 32.45222, 37.20556, 40.86639, 42.93972, 
    18.43083, 25.91556, 27.77944, 32.12361, 32.84444, 39.56861, 40.77389, 
    42.38139, 44.90833, 44.84722, 44.07778, 47.46028, 47.9375, 41.6125, 
    7.08694, 9.48333, 8.73333, 82.5, 50.23, 53.3, 51.48, 53.98, 63.76, 74.72, 
    60.04, 68.32, 60.73, 65.28, 51.28, 12.2, 49.97, 43.94, 80, 69.1, 24.3, 
    50.69, 53.55, 17.5, 32.85, 17.93333, 52.73, 33.26, 34.93, 13.55, 16.733, 
    -9.817 ;

 staLon = -64.68333, -77.46667, -156.8025, -117.9, -120.57, -120.5667, 
    158.2167, -122.6, -165.4403, -170.2167, -162.7233, -156.6683, -152.4833, 
    -159.35, 134.4833, -86.78361, -162.6333, -161.8442, -155.6167, -147.8772, 
    -149.9864, -139.6719, -131.5781, -155.0667, 151.8364, -82.40194, 
    -108.4767, -100.7611, -170.7167, -52.75, -96, -80.38389, -90.08028, 
    -76.87917, -79.95, -86.55, -75.48333, -83.82111, -73.8, -80.21806, 
    -83.47167, -68.01667, -70.25787, -69.96667, -89.33861, -89.83056, 
    -97.29722, -100.9167, -102.1889, -92.25861, -97.46083, -101.7083, 
    -106.6833, -106.6219, -111.8203, -116.0217, -93.40194, -99.96889, 
    -104.8694, -108.5333, -122.2206, -96.36611, -100.7006, -115.7417, 
    -88.11083, -98.41389, -116.2264, -93.39694, -106.625, -117.6258, 
    144.7975, -81.25, -66.08, -75.97, -58.55, -68.42, -78.12, -77.46667, 
    -81.75, -81.70167, -80.03333, -84.35056, -84.56722, -93.21639, -93.8425, 
    -80.41417, -72.85139, -78.73611, -65.99167, -97.41972, -97.505, 
    -110.9425, -117.1233, -119.7964, -111.9544, -122.8778, -84.71944, 
    -93.56444, -103.2167, -111.3842, -124.555, -90.58222, 171.3875, 138.0833, 
    167.7333, -62.33, -66.27, -60.37, -90.2, -101.1, -68.55, -94.95, -111.93, 
    -133.53, -135.07, -126.8, -80.65, -68.96667, -119.38, -60.02, -85.93, 
    -105.12, 153.967, -127.37, -114.1, -88.33333, -114.4, -76.78333, 174.1, 
    -119.45, -117.9, 144.833, -169.51, -139.01 ;

 staElev = 6, 2, 12, 705, 100, 112, 39, 382, 5, 10, 30, 15, 4, 32, 30, 174, 
    5, 36, 103, 135, 50, 12, 37, 10, 3, 13, 1700, 505, 5, 140, 49, 5, 91, 11, 
    277, 180, 13, 323, 86, 360, 329, 191, 125, 16, 178, 10, 198, 314, 873, 
    172, 357, 1094, 1257, 1615, 2180, 1007, 390, 790, 1611, 1475, 6, 350, 
    847, 1607, 214, 397, 871, 361, 692, 728, 90, 7, 43, 170, 61, 36, 7, 85, 
    2, 11, 15, 18, 246, 5, 85, 0, 20, 218, 3, 7, 14, 787, 134, 1516, 1288, 
    397, 1465, 288, 1027, 1132, 56, 229, 3, 14, 8, 66, 53, 36, 373, 273, 21, 
    40, 203, 68, 700, 60, 10, 62, 429, 4, 10, 25, 8, 17, 766, 5, 98, 3, 39, 
    153, 705, 111, 3, 52 ;

 synTime = 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 1085054400, 
    1085054400, 1085054400, 1085054400, 1085054400, 1085058000, 1085058000, 
    1085054400, 1085054400, 1085054400 ;

 numMand = 0, 12, 12, 0, 12, 0, 12, 12, 12, 12, 12, 12, 12, 12, 12, 0, 12, 
    12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 
    12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 
    12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 
    12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 
    12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 
    12, 12, 12, 12, 12, 12, 12, _, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 
    12, 12, 12, 12, 12, 12, 0, 0, 12 ;

 numSigT = _, 14, 10, _, 35, _, _, 28, 23, 13, 16, 21, 21, 27, 23, _, 21, 24, 
    24, 27, 23, 15, 14, 34, 13, 26, 19, 31, 34, 20, 31, 20, 32, 26, 21, 27, 
    20, 16, 19, 20, 21, 16, 21, 13, 18, 30, 13, 14, 13, 17, 18, 22, 15, 18, 
    19, 10, 20, 14, 18, 16, 21, 19, 24, 16, 20, 22, 16, 24, 20, 15, 27, 25, 
    23, 24, 23, 17, 25, 25, 28, 20, 19, 18, 20, 22, 20, 18, 20, 20, 28, 13, 
    18, 16, 21, 14, 25, 27, 28, 28, 18, 19, 20, 17, 22, 31, 11, 25, 28, 23, 
    28, 26, 21, 27, 29, 23, 27, 18, 18, 22, 26, 22, 20, _, 17, 27, 21, 30, 
    19, 32, 22, 17, 12, _, _, 17 ;

 numSigW = _, 26, 23, _, 30, _, 26, 22, 20, 20, 23, 21, 22, 27, 23, _, 21, 
    20, 21, 22, 23, 22, 23, 24, 27, 22, 18, 24, 25, 26, 26, 24, 30, 24, 22, 
    28, 25, 24, 27, 24, 27, 20, 24, 22, 22, 27, 23, 21, 23, 22, 25, 22, 24, 
    23, 15, 22, 25, 23, 16, 19, 23, 24, 21, 15, 22, 24, 21, 24, 22, 22, 25, 
    30, 23, 25, 28, 26, 26, 23, 20, 25, 30, 16, 24, 17, 25, 28, 25, 21, 26, 
    20, 23, 22, 21, 19, 18, 20, 24, 24, 16, 22, 27, 22, 23, 27, 17, 22, 26, 
    25, 23, 23, 30, 23, 18, 24, 23, 28, 26, 10, 30, 30, 30, 19, _, 27, 30, 
    30, 17, 17, 23, 6, 19, _, _, _ ;

 numMwnd = 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 
    1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 
    0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 
    1, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, _, 0, 1, 0, 
    0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0 ;

 numTrop = 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 2, 1, 1, 1, 1, 2, _, 1, 2, 1, 
    1, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0 ;

 relTime = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 sondTyp = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 prMan =
  0, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 
    10000, 0, _, _, _, _, _, _, _, _, _,
  1021, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1029, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  0, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 
    10000, -99999, _, _, _, _, _, _, _, _, _,
  1005, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, -99999, _, _, 
    _, _, _, _, _, _, _,
  0, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 
    10000, -99999, _, _, _, _, _, _, _, _, _,
  1007, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  979, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1034, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1025, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1024, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1031, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1031, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1011, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1008, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  0, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 
    10000, 0, _, _, _, _, _, _, _, _, _,
  1032, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1028, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1019, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1015, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1025, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1025, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1015, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1014, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1011, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1021, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  831, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  960, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1012, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1004, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1010, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1021, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1012, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1021, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  990, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1000, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1022, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  981, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1014, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  979, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  977, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1001, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1010, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1024, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  993, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1021, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  995, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  979, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  917, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  999, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  974, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  893, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  875, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  839, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  784, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  896, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  972, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  922, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  840, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  849, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1015, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  970, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  919, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  838, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  985, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  970, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  915, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  969, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  937, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  931, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1004, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1011, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1025, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  997, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1017, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1001, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  997, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1013, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1020, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1022, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1021, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1017, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  995, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1021, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1011, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  949, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1023, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  993, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1017, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1016, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1016, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  924, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1000, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  847, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  866, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  969, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  959, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  976, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  901, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  888, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1012, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  985, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1011, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1009, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1010, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1016, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1017, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1015, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  966, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  992, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1006, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1015, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1004, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1019, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1017, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1004, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1008, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  961, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1025, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1020, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1022, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1015, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1017, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  931, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1016, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  992, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  1015, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1016, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  1016, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _,
  930, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, _, 
    _, _, _, _, _,
  0, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 
    10000, 0, _, _, _, _, _, _, _, _, _,
  0, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 
    10000, 0, _, _, _, _, _, _, _, _, _,
  1007, 1000, 925, 850, 700, 500, 400, 300, 250, 200, 150, 100, _, _, _, _, 
    _, _, _, _, _, _ ;

 htMan =
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 2.003573, _, _, _, _, _, _, _, _, _,
  2, -99999, -99999, 1577, 3185, 5870, 7550, 9600, 10830, 12280, 14070, 
    16530, _, _, _, _, _, _, _, _, _, _,
  12, 241, 867, 1533, 3017, 5470, 7010, 8910, 10110, 11610, 13540, 16230, _, 
    _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 2.003573, _, _, _, _, _, _, _, _, _,
  100, 141, 786, 1490, 3074, 5680, 7310, 9300, 10500, 11970, 13820, 16400, 
    2.003573, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 2.003573, _, _, _, _, _, _, _, _, _,
  39, 99, 785, 1518, 3164, 5890, 7610, 9720, 10990, 12470, 14260, 16620, _, 
    _, _, _, _, _, _, _, _, _,
  382, 209, 850, 1533, 3065, 5590, 7160, 9080, 10250, 11700, 13590, 16230, _, 
    _, _, _, _, _, _, _, _, _,
  5, 271, 894, 1562, 3058, 5580, 7150, 9100, 10280, 11730, 13620, 16270, _, 
    _, _, _, _, _, _, _, _, _,
  10, 212, 845, 1524, 3069, 5670, 7310, 9300, 10500, 11910, 13700, 16300, _, 
    _, _, _, _, _, _, _, _, _,
  30, 222, 854, 1548, 3122, 5740, 7380, 9390, 10610, 12020, 13790, 16360, _, 
    _, _, _, _, _, _, _, _, _,
  15, 264, 904, 1589, 3153, 5760, 7400, 9400, 10620, 12040, 13800, 16370, _, 
    _, _, _, _, _, _, _, _, _,
  4, 258, 900, 1593, 3164, 5790, 7430, 9420, 10640, 12060, 13820, 16380, _, 
    _, _, _, _, _, _, _, _, _,
  32, 124, 803, 1528, 3151, 5850, 7550, 9620, 10860, 12320, 14110, 16510, _, 
    _, _, _, _, _, _, _, _, _,
  30, 97, 784, 1516, 3161, 5890, 7610, 9720, 10980, 12460, 14260, 16620, _, 
    _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 2.003573, _, _, _, _, _, _, _, _, _,
  5, 261, 884, 1549, 3036, 5520, 7080, 9000, 10190, 11670, 13580, 16260, _, 
    _, _, _, _, _, _, _, _, _,
  36, 265, 903, 1583, 3121, 5700, 7330, 9320, 10520, 11940, 13730, 16330, _, 
    _, _, _, _, _, _, _, _, _,
  103, 260, 901, 1582, 3100, 5660, 7270, 9250, 10440, 11850, 13680, 16300, _, 
    _, _, _, _, _, _, _, _, _,
  135, 258, 901, 1584, 3095, 5600, 7190, 9130, 10320, 11760, 13640, 16280, _, 
    _, _, _, _, _, _, _, _, _,
  50, 252, 897, 1583, 3134, 5720, 7360, 9340, 10540, 11950, 13750, 16340, _, 
    _, _, _, _, _, _, _, _, _,
  12, 215, 856, 1555, 3126, 5720, 7350, 9330, 10530, 11930, 13730, 16320, _, 
    _, _, _, _, _, _, _, _, _,
  37, 164, 821, 1529, 3111, 5720, 7360, 9350, 10550, 11960, 13740, 16320, _, 
    _, _, _, _, _, _, _, _, _,
  10, 134, 813, 1537, 3172, 5870, 7570, 9640, 10890, 12340, 14130, 16530, _, 
    _, _, _, _, _, _, _, _, _,
  3, 96, 781, 1512, 3155, 5890, 7600, 9700, 10970, 12440, 14230, 16570, _, _, 
    _, _, _, _, _, _, _, _,
  13, 192, 866, 1587, 3196, 5880, 7560, 9610, 10830, 12260, 14000, 16470, _, 
    _, _, _, _, _, _, _, _, _,
  1700, 98, 778, 1504, 3093, 5720, 7370, 9370, 10580, 11990, 13800, 16350, _, 
    _, _, _, _, _, _, _, _, _,
  505, 154, 813, 1508, 3076, 5680, 7330, 9340, 10550, 11980, 13780, 16350, _, 
    _, _, _, _, _, _, _, _, _,
  5, 108, 796, 1529, 3173, 5890, 7590, 9680, 10940, 12400, 14180, 16550, _, 
    _, _, _, _, _, _, _, _, _,
  140, 174, 805, 1483, 3007, 5560, 7170, 9140, 10330, 11780, 13650, 16260, _, 
    _, _, _, _, _, _, _, _, _,
  49, 130, 732, 1374, 2844, 5300, 6830, 8700, -99999, 11410, 13360, 16080, _, 
    _, _, _, _, _, _, _, _, _,
  5, 185, 859, 1579, 3191, 5870, 7550, 9590, 10810, 12250, 14030, 16480, _, 
    _, _, _, _, _, _, _, _, _,
  91, 192, 868, 1591, 3213, 5890, 7570, 9640, 10880, 12320, 14070, 16510, _, 
    _, _, _, _, _, _, _, _, _,
  11, 194, 869, 1591, 3201, 5870, 7550, 9600, 10820, 12250, 13980, 16430, _, 
    _, _, _, _, _, _, _, _, _,
  277, 188, 863, 1587, 3200, 5870, 7550, 9600, 10820, 12250, 13990, 16420, _, 
    _, _, _, _, _, _, _, _, _,
  180, 180, 860, 1583, 3205, 5880, 7570, 9630, 10860, 12300, 14060, 16490, _, 
    _, _, _, _, _, _, _, _, _,
  13, 194, 856, 1567, 3174, 5850, 7530, 9560, 10780, 12200, 13950, 16410, _, 
    _, _, _, _, _, _, _, _, _,
  323, 156, 832, 1556, 3171, 5860, 7540, 9580, 10810, 12240, 13990, 16410, _, 
    _, _, _, _, _, _, _, _, _,
  86, 204, 859, 1562, 3148, 5800, 7460, 9480, 10680, 12100, 13860, 16370, _, 
    _, _, _, _, _, _, _, _, _,
  360, 173, 841, 1559, 3165, 5830, 7520, 9560, 10790, 12220, 13980, 16430, _, 
    _, _, _, _, _, _, _, _, _,
  329, 129, 796, 1517, 3133, 5800, 7470, 9510, 10740, 12160, 13910, 16380, _, 
    _, _, _, _, _, _, _, _, _,
  191, 199, 850, 1548, 3108, 5700, 7320, 9320, 10520, 11930, 13730, 16290, _, 
    _, _, _, _, _, _, _, _, _,
  125, 210, 868, 1568, 3137, 5750, 7400, 9410, 10600, 12020, 13780, 16300, _, 
    _, _, _, _, _, _, _, _, _,
  16, 214, 869, 1567, 3146, 5780, 7440, 9450, 10650, 12050, 13830, 16350, _, 
    _, _, _, _, _, _, _, _, _,
  178, 118, 795, 1523, 3155, 5850, 7540, 9580, 10810, 12240, 13990, 16410, _, 
    _, _, _, _, _, _, _, _, _,
  10, 190, 866, 1588, 3210, 5880, 7560, 9620, 10850, 12280, 14040, 16480, _, 
    _, _, _, _, _, _, _, _, _,
  198, 153, 829, 1556, 3191, 5900, 7590, 9640, 10870, 12310, 14080, 16500, _, 
    _, _, _, _, _, _, _, _, _,
  314, 130, 811, 1535, 3165, 5890, 7580, 9650, 10900, 12350, 14140, 16570, _, 
    _, _, _, _, _, _, _, _, _,
  873, 94, 792, 1521, 3167, 5880, 7570, 9620, 10860, 12300, 14070, 16510, _, 
    _, _, _, _, _, _, _, _, _,
  172, 165, 841, 1569, 3213, 5900, 7570, 9630, 10860, 12310, 14050, 16470, _, 
    _, _, _, _, _, _, _, _, _,
  357, 120, 801, 1534, 3194, 5890, 7570, 9610, 10840, 12290, 14030, 16460, _, 
    _, _, _, _, _, _, _, _, _,
  1094, 86, 782, 1516, 3174, 5870, 7560, 9610, 10840, 12270, 14030, 16480, _, 
    _, _, _, _, _, _, _, _, _,
  1257, 47, 753, 1504, 3163, 5860, 7530, 9600, 10830, 12270, 14050, 16500, _, 
    _, _, _, _, _, _, _, _, _,
  1615, 41, 745, 1498, 3150, 5840, 7510, 9560, 10790, 12230, 14000, 16500, _, 
    _, _, _, _, _, _, _, _, _,
  2180, 96, 773, 1496, 3109, 5780, 7450, 9490, 10700, 12130, 13900, 16450, _, 
    _, _, _, _, _, _, _, _, _,
  1007, 37, 727, 1454, 3063, 5700, 7340, 9350, 10560, 11990, 13840, 16420, _, 
    _, _, _, _, _, _, _, _, _,
  390, 140, 817, 1545, 3205, 5890, 7570, 9620, 10840, 12280, 14030, 16450, _, 
    _, _, _, _, _, _, _, _, _,
  790, 62, 758, 1501, 3166, 5870, 7550, 9600, 10830, 12260, 14010, 16470, _, 
    _, _, _, _, _, _, _, _, _,
  1611, 75, 770, 1512, 3135, 5800, 7460, 9500, 10720, 12150, 13910, 16410, _, 
    _, _, _, _, _, _, _, _, _,
  1475, 20, 718, 1463, 3108, 5770, 7440, 9470, 10680, 12110, 13890, 16420, _, 
    _, _, _, _, _, _, _, _, _,
  6, 134, 779, 1479, 3054, 5650, 7260, 9220, 10420, 11870, 13750, 16350, _, 
    _, _, _, _, _, _, _, _, _,
  350, 87, 762, 1494, 3141, 5830, 7510, 9540, 10760, 12200, 13960, 16420, _, 
    _, _, _, _, _, _, _, _, _,
  847, 110, 791, 1502, 3133, 5820, 7480, 9520, 10740, 12180, 13920, 16420, _, 
    _, _, _, _, _, _, _, _, _,
  1607, 73, 747, 1467, 3064, 5670, 7290, 9270, 10460, 11900, 13760, 16350, _, 
    _, _, _, _, _, _, _, _, _,
  214, 84, 751, 1472, 3091, 5750, 7430, 9480, 10720, 12160, 13910, 16400, _, 
    _, _, _, _, _, _, _, _, _,
  397, 131, 790, 1487, 3072, 5720, 7380, 9400, 10620, 12050, 13820, 16350, _, 
    _, _, _, _, _, _, _, _, _,
  871, 110, 775, 1479, 3056, 5650, 7260, 9210, 10400, 11850, 13710, 16300, _, 
    _, _, _, _, _, _, _, _, _,
  361, 90, 742, 1435, 3002, 5610, 7260, 9260, 10470, 11900, 13720, 16300, _, 
    _, _, _, _, _, _, _, _, _,
  692, 142, 801, 1512, 3090, 5670, 7290, 9260, 10460, 11870, 13720, 16310, _, 
    _, _, _, _, _, _, _, _, _,
  728, 120, 782, 1485, 3063, 5650, 7270, 9230, 10400, 11820, 13680, 16270, _, 
    _, _, _, _, _, _, _, _, _,
  90, 106, 793, 1527, 3171, 5880, 7590, 9670, 10930, 12400, 14200, 16590, _, 
    _, _, _, _, _, _, _, _, _,
  7, 91, 702, 1356, 2834, 5290, 6840, 8740, -99999, 11430, 13360, 16090, _, 
    _, _, _, _, _, _, _, _, _,
  43, 215, 868, 1567, 3124, 5730, 7370, 9370, 10560, 11960, 13770, 16320, _, 
    _, _, _, _, _, _, _, _, _,
  170, 163, 819, 1521, 3106, 5720, 7380, 9410, 10620, 12040, 13810, 16320, _, 
    _, _, _, _, _, _, _, _, _,
  61, 195, 829, 1508, 3031, 5570, 7160, 9110, 10290, 11730, 13610, 16230, _, 
    _, _, _, _, _, _, _, _, _,
  36, 71, 697, 1373, 2906, 5450, 7050, 8980, 10150, 11580, 13460, 16130, _, 
    _, _, _, _, _, _, _, _, _,
  7, 1, 608, 1276, 2799, 5340, 6930, 8880, 10060, 11510, 13420, 16110, _, _, 
    _, _, _, _, _, _, _, _,
  85, 198, 862, 1574, 3178, 5850, 7530, 9570, 10790, 12210, 13960, 16420, _, 
    _, _, _, _, _, _, _, _, _,
  2, 178, 854, 1574, 3191, 5880, 7560, 9600, 10840, 12280, 14070, 16530, _, 
    _, _, _, _, _, _, _, _, _,
  11, 199, 873, 1592, 3201, 5880, 7560, 9610, 10830, 12260, 14000, 16440, _, 
    _, _, _, _, _, _, _, _, _,
  15, 199, 874, 1595, 3208, 5880, 7570, 9610, 10840, 12270, 14020, 16460, _, 
    _, _, _, _, _, _, _, _, _,
  18, 195, 870, 1593, 3206, 5870, 7550, 9600, 10830, 12260, 14000, 16440, _, 
    _, _, _, _, _, _, _, _, _,
  246, 200, 874, 1596, 3210, 5880, 7560, 9620, 10850, 12280, 14020, 16440, _, 
    _, _, _, _, _, _, _, _, _,
  5, 183, 858, 1581, 3205, 5880, -99999, -99999, -99999, -99999, -99999, 
    -99999, _, _, _, _, _, _, _, _, _, _,
  85, 179, 851, 1575, 3203, 5890, 7570, 9630, 10860, 12300, 14050, 16470, _, 
    _, _, _, _, _, _, _, _, _,
  0, 191, 862, 1584, 3198, 5870, 7560, 9610, 10830, 12260, 14000, 16430, _, 
    _, _, _, _, _, _, _, _, _,
  20, 214, 869, 1569, 3157, 5810, 7480, 9490, 10690, 12100, 13860, 16360, _, 
    _, _, _, _, _, _, _, _, _,
  218, 161, 825, 1538, 3135, 5790, 7470, 9500, 10720, 12130, 13890, 16360, _, 
    _, _, _, _, _, _, _, _, _,
  3, 153, 833, 1556, 3182, 5880, 7590, 9690, 10950, 12420, 14210, 16570, _, 
    _, _, _, _, _, _, _, _, _,
  7, 147, 826, 1549, 3177, 5880, 7580, 9660, 10900, 12360, 14150, 16570, _, 
    _, _, _, _, _, _, _, _, _,
  14, 152, 830, 1553, 3178, 5890, 7590, 9660, 10900, 12360, 14140, 16560, _, 
    _, _, _, _, _, _, _, _, _,
  787, 78, 775, 1507, 3143, 5820, 7500, 9550, 10780, 12220, 14010, 16490, _, 
    _, _, _, _, _, _, _, _, _,
  134, 131, 787, 1488, 3086, 5740, 7410, 9440, 10660, 12090, 13880, 16440, _, 
    _, _, _, _, _, _, _, _, _,
  1516, 99, 768, 1482, 3062, 5650, 7250, 9200, 10400, 11850, 13730, 16330, _, 
    _, _, _, _, _, _, _, _, _,
  1288, 37, 720, 1447, 3068, 5700, 7350, 9350, 10560, 11970, 13780, 16350, _, 
    _, _, _, _, _, _, _, _, _,
  397, 131, 786, 1487, 3060, 5640, 7260, 9210, 10380, 11830, 13700, 16300, _, 
    _, _, _, _, _, _, _, _, _,
  1465, 85, 747, 1466, 3073, 5740, 7410, 9460, 10680, 12100, 13850, 16350, _, 
    _, _, _, _, _, _, _, _, _,
  288, 84, 752, 1471, 3081, 5750, 7410, 9450, 10670, 12100, 13860, 16370, _, 
    _, _, _, _, _, _, _, _, _,
  1027, 131, 805, 1515, 3105, 5740, 7390, 9410, 10620, 12050, 13820, 16350, 
    _, _, _, _, _, _, _, _, _, _,
  1132, 136, 791, 1493, 3074, 5660, 7280, 9240, 10430, 11850, 13690, 16290, 
    _, _, _, _, _, _, _, _, _, _,
  56, 159, 802, 1502, 3090, 5680, 7300, 9280, 10470, 11870, 13710, 16280, _, 
    _, _, _, _, _, _, _, _, _,
  229, 94, 773, 1503, 3138, 5830, 7510, 9560, 10780, 12210, 13970, 16390, _, 
    _, _, _, _, _, _, _, _, _,
  3, 99, 785, 1516, 3160, 5890, 7610, 9710, 10980, 12460, 14260, 16610, _, _, 
    _, _, _, _, _, _, _, _,
  14, 94, 780, 1513, 3157, 5880, 7590, 9700, 10960, 12440, 14230, 16580, _, 
    _, _, _, _, _, _, _, _, _,
  8, 95, 786, 1522, 3171, 5890, 7610, 9720, 10990, 12480, 14270, 16620, _, _, 
    _, _, _, _, _, _, _, _,
  66, 189, 792, 1459, 2967, 5440, 7000, 8910, 10080, 11550, 13470, 16180, _, 
    _, _, _, _, _, _, _, _, _,
  53, 189, 829, 1514, 3060, 5630, 7230, 9210, 10390, 11790, 13620, 16220, _, 
    _, _, _, _, _, _, _, _, _,
  36, 160, 787, 1454, 2965, 5480, 7060, 8980, 10160, 11600, 13500, 16150, _, 
    _, _, _, _, _, _, _, _, _,
  373, 109, 728, 1393, 2932, 5500, 7120, 9090, 10280, 11730, 13610, 16220, _, 
    _, _, _, _, _, _, _, _, _,
  273, 208, 817, 1476, 2976, 5490, 7080, 9010, 10190, 11650, 13540, 16190, _, 
    _, _, _, _, _, _, _, _, _,
  21, 69, 686, 1345, 2836, 5330, 6890, 8790, -99999, 11460, 13380, 16100, _, 
    _, _, _, _, _, _, _, _, _,
  40, 158, 763, 1415, 2910, 5380, 6940, 8850, 10030, 11520, 13440, 16150, _, 
    _, _, _, _, _, _, _, _, _,
  203, 233, 843, 1497, 2988, 5470, 7030, 8930, 10110, 11570, 13480, 16150, _, 
    _, _, _, _, _, _, _, _, _,
  68, 248, 870, 1538, 3036, 5500, 7040, 8940, 10140, 11620, 13550, 16230, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  60, 233, 856, 1526, 3032, 5510, 7050, 8950, 10140, 11630, 13540, 16220, _, 
    _, _, _, _, _, _, _, _, _,
  10, 42, 695, 1393, 2945, 5540, 7170, 9160, 10350, 11790, 13630, 16210, _, 
    _, _, _, _, _, _, _, _, _,
  62, 124, 812, -99999, -99999, 5880, -99999, 9710, 10980, 12460, 14250, 
    16600, _, _, _, _, _, _, _, _, _, _,
  429, 123, 780, 1488, 3074, 5660, 7270, 9230, 10410, 11820, 13680, 16270, _, 
    _, _, _, _, _, _, _, _, _,
  4, 206, 848, 1535, 3091, 5680, 7310, 9300, 10500, 11920, 13730, 16290, _, 
    _, _, _, _, _, _, _, _, _,
  10, 167, 781, 1449, 2960, 5460, 7020, 8930, 10110, 11590, 13500, 16190, _, 
    _, _, _, _, _, _, _, _, _,
  25, 193, 778, 1423, 2912, 5390, 6940, 8840, 10020, 11490, 13430, 16150, _, 
    _, _, _, _, _, _, _, _, _,
  8, 135, 813, 1536, 3177, 5910, 7620, 9710, 10980, 12450, 14240, 16620, _, 
    _, _, _, _, _, _, _, _, _,
  17, 158, 802, 1510, 3097, 5710, 7350, 9340, 10530, 11940, 13740, 16310, _, 
    _, _, _, _, _, _, _, _, _,
  766, 176, 822, 1509, 3052, 5610, 7210, 9150, 10310, 11730, 13600, 16220, _, 
    _, _, _, _, _, _, _, _, _,
  5, 140, 832, 1554, 3186, 5900, 7610, 9710, 10990, 12460, 14250, 16620, _, 
    _, _, _, _, _, _, _, _, _,
  98, 63, 741, 1467, 3095, 5760, 7430, 9470, 10700, 12130, -99999, -99999, _, 
    _, _, _, _, _, _, _, _, _,
  3, 132, -99999, 1544, 3173, -99999, -99999, -99999, -99999, 12420, 14210, 
    16540, _, _, _, _, _, _, _, _, _, _,
  39, 157, 791, 1476, 3009, 5550, 7150, 9080, 10250, 11690, -99999, -99999, 
    _, _, _, _, _, _, _, _, _, _,
  153, 149, 796, 1503, 3096, 5720, 7370, 9390, 10610, 12050, -99999, -99999, 
    _, _, _, _, _, _, _, _, _, _,
  705, 105, -99999, 1471, 3066, 5690, 7330, 9330, 10540, 11990, 13820, 16400, 
    _, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 2.003573, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 2.003573, _, _, _, _, _, _, _, _, _,
  52, 108, 790, 1517, 3152, 5870, 7590, 9690, 10940, 12410, 14190, 16570, _, 
    _, _, _, _, _, _, _, _, _ ;

 tpMan =
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 0, _, _, _, _, _, _, _, _, _,
  296.1, -99999, -99999, 286.1, 278.5, 263.8, 250.6, 235.4, 226.2, 217.2, 
    208.6, 205.4, _, _, _, _, _, _, _, _, _, _,
  272.6, 275.9, 271, 266.6, 256, 241.8, 231.2, 222.8, 227.2, 229.2, 229.4, 
    224.2, _, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 0, _, _, _, _, _, _, _, _, _,
  283.9, -99999, 280.5, 283.5, 274.9, 255.4, 243.8, 228.8, 224.8, 221.8, 
    218.8, 216, 0, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 0, _, _, _, _, _, _, _, _, _,
  297.7, 298.7, 295.3, 291.7, 283.5, 268.4, 257.6, 242.4, 232.2, 220, 206.8, 
    194, _, _, _, _, _, _, _, _, _, _,
  280.9, -99999, 277.5, 272.8, 263.8, 247.8, 235.6, 221, 218.6, 222.8, 224.4, 
    220.6, _, _, _, _, _, _, _, _, _, _,
  274.1, 273.3, 271.2, 266.6, 261, 247.8, 237, 224, 220.6, 224.4, 224.4, 221, 
    _, _, _, _, _, _, _, _, _, _,
  277.5, 277.1, 275.3, 272.4, 270, 256.6, 244.2, 229, 220.2, 210.6, 216.2, 
    219, _, _, _, _, _, _, _, _, _, _,
  278.7, 277.7, 275.7, 280.3, 272.2, 257, 246.6, 231, 222.2, 211.4, 212.8, 
    216.8, _, _, _, _, _, _, _, _, _, _,
  279.5, 279.7, 277.9, 276.3, 272.6, 257, 244.8, 231, 223, 211.6, 212.8, 
    217.8, _, _, _, _, _, _, _, _, _, _,
  279.7, 281.3, 280.5, 278.1, 273.1, 257, 244.6, 231, 222.8, 211.2, 213.8, 
    216.2, _, _, _, _, _, _, _, _, _, _,
  298.1, 297.3, 292.7, 288.5, 279.7, 266.2, 254.6, 237.4, 228.4, 217.6, 
    207.6, 200, _, _, _, _, _, _, _, _, _, _,
  300.3, 300.1, 295.5, 291.9, 283.9, 267.6, 258.2, 241.6, 232.4, 220.4, 206, 
    193.2, _, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 0, _, _, _, _, _, _, _, _, _,
  274.7, 274.3, 270.2, 265.2, 258.4, 243.6, 234.6, 223.8, 224.4, 226.6, 
    226.2, 223.4, _, _, _, _, _, _, _, _, _, _,
  278.1, 281.5, 276.3, 271, 267.6, 254.4, 243.6, 229.4, 222.4, 211.8, 216.8, 
    220.2, _, _, _, _, _, _, _, _, _, _,
  278.1, 281.3, 277.5, 271.4, 264, 251.6, 241.8, 227.8, 220.6, 212.8, 218.6, 
    220.2, _, _, _, _, _, _, _, _, _, _,
  279.1, 280.9, 278.7, 271.8, 260, 248.4, 237.2, 223.4, 221, 221.4, 223.2, 
    221.8, _, _, _, _, _, _, _, _, _, _,
  280.1, 282.7, 279.3, 274.3, 270, 255.4, 243.8, 228.8, 221.2, 209.8, 217.6, 
    220.2, _, _, _, _, _, _, _, _, _, _,
  278.1, 278.9, 280.9, 281.3, 271, 254.8, 243.2, 227.6, 220, 209.2, 218, 
    218.2, _, _, _, _, _, _, _, _, _, _,
  284.1, 286.7, 287.5, 282.9, 273.1, 256.6, 244.2, 228.8, 220.2, 211, 216, 
    215.8, _, _, _, _, _, _, _, _, _, _,
  295.9, 297.1, 292.5, 289.5, 281.1, 265, 254.4, 238, 227.6, 216.8, 207.8, 
    200.8, _, _, _, _, _, _, _, _, _, _,
  300.7, 300.3, 294.7, 290.5, 283.9, 267.4, 256.6, 241.8, 232.2, 219, 204, 
    194.6, _, _, _, _, _, _, _, _, _, _,
  293.5, 294.9, 291.9, 286.7, 278.5, 263, 251.4, 234.8, 224.2, 212.4, 208, 
    204.4, _, _, _, _, _, _, _, _, _, _,
  281.3, -99999, -99999, -99999, 273.5, 257.4, 245.6, 230.8, 221.4, 213, 
    215.2, 214.2, _, _, _, _, _, _, _, _, _, _,
  283.1, -99999, 281.5, 277.5, 272.8, 256, 246.2, 231, 223.2, 214, 214.4, 
    217.6, _, _, _, _, _, _, _, _, _, _,
  299.7, 300.1, 296.1, 291.9, 283.5, 266.2, 255, 240.6, 230.8, 217.6, 205.2, 
    198.6, _, _, _, _, _, _, _, _, _, _,
  279.1, 278.3, 275.1, 270.8, 265.6, 252.2, 240.4, 226.4, 221.6, 219.6, 
    220.6, 219.6, _, _, _, _, _, _, _, _, _, _,
  263.4, 262.8, 262.4, 256.6, 256.6, 240.6, 228, 220.8, 228.6, 231.2, 230.2, 
    228.6, _, _, _, _, _, _, _, _, _, _,
  295.5, 296.1, 290.7, 287.5, 279.7, 263.2, 250.4, 234.2, 224.8, 214.6, 209, 
    205.6, _, _, _, _, _, _, _, _, _, _,
  291.9, 293.3, 292.5, 289.1, 280.1, 262.4, 252.4, 237, 226.8, 214.4, 203.2, 
    205.6, _, _, _, _, _, _, _, _, _, _,
  294.7, 294.3, 292.1, 287.3, 278.3, 262.4, 252, 234, 223.8, 212, 205.4, 
    209.6, _, _, _, _, _, _, _, _, _, _,
  291.3, -99999, 293.3, 287.9, 277.9, 263.2, 252.2, 234.2, 224.2, 213, 201.4, 
    206.4, _, _, _, _, _, _, _, _, _, _,
  292.1, 292.1, 292.5, 287.9, 279.9, 263, 252.2, 236.2, 225.4, 215.4, 202.6, 
    208, _, _, _, _, _, _, _, _, _, _,
  289.7, 288.5, 286.9, 284.1, 278.3, 262.6, 249.8, 232.6, 222.4, 212.4, 
    208.2, 208, _, _, _, _, _, _, _, _, _, _,
  293.1, -99999, 292.5, 287.7, 278.3, 264.6, 250.6, 234, 225.2, 213.4, 202.4, 
    206.4, _, _, _, _, _, _, _, _, _, _,
  281.9, 282.1, 285.9, 280.1, 274.5, 260.4, 247.8, 231, 220.8, 212, 210.6, 
    211.6, _, _, _, _, _, _, _, _, _, _,
  289.1, -99999, 290.1, 286.3, 276.5, 263.2, 251.2, 234.6, 225, 213.2, 204.4, 
    210, _, _, _, _, _, _, _, _, _, _,
  287.3, -99999, 290.9, 286.5, 279.1, 260, 250, 234.8, 224.4, 211.8, 207.6, 
    210.2, _, _, _, _, _, _, _, _, _, _,
  279.7, 279.7, 284.5, 278.3, 270.2, 253.4, 243, 229, 220.6, 212.2, 215.6, 
    217.2, _, _, _, _, _, _, _, _, _, _,
  284.5, 286.9, 285.1, 278.9, 272, 258.2, 246.6, 229.4, 221.2, 210.4, 210.6, 
    212, _, _, _, _, _, _, _, _, _, _,
  285.5, 288.3, 284.1, 279.1, 273.7, 261.8, 247.4, 230, 219.4, 210, 210.4, 
    212.2, _, _, _, _, _, _, _, _, _, _,
  293.9, -99999, 293.7, 289.5, 284.1, 264, 250, 234.4, 224.6, 214.4, 201.8, 
    207.6, _, _, _, _, _, _, _, _, _, _,
  291.3, 295.5, 292.1, 289.1, 278.9, 262.2, 252, 235.6, 225.6, 214.4, 203, 
    205, _, _, _, _, _, _, _, _, _, _,
  295.3, -99999, 292.9, 290.3, 283.7, 265.4, 252.8, 235.4, 225.8, 215.4, 
    204.4, 203.8, _, _, _, _, _, _, _, _, _, _,
  295.9, -99999, 292.1, 289.7, 285.9, 266.2, 252.8, 239.2, 228.2, 216.8, 
    207.4, 202, _, _, _, _, _, _, _, _, _, _,
  293.3, -99999, -99999, 288.9, 285.5, 264.2, 252.4, 237.2, 226.6, 215.4, 
    206.6, 203.6, _, _, _, _, _, _, _, _, _, _,
  293.7, -99999, 294.1, 290.1, 283.1, 261, 251.4, 236.2, 226, 214.4, 200.6, 
    205, _, _, _, _, _, _, _, _, _, _,
  294.3, -99999, 294.9, 295.5, 284.9, 263.8, 250.8, 233.6, 226.6, 214.8, 
    202.8, 203.6, _, _, _, _, _, _, _, _, _, _,
  290.7, -99999, -99999, 291.3, 284.9, 263.6, 250.6, 235.4, 225.6, 213.8, 
    205, 205.2, _, _, _, _, _, _, _, _, _, _,
  295.1, -99999, -99999, 296.3, 284.3, 262, 253.6, 236.2, 225.6, 215.8, 207, 
    202.4, _, _, _, _, _, _, _, _, _, _,
  293.3, -99999, -99999, -99999, 283.5, 260.4, 251.8, 235.6, 226, 214.4, 
    210.2, 206.6, _, _, _, _, _, _, _, _, _, _,
  273.5, -99999, -99999, -99999, 278.1, 262.4, 250.2, 233, 223.4, 211.6, 
    214.6, 209.4, _, _, _, _, _, _, _, _, _, _,
  291.1, -99999, -99999, 288.3, 276.3, 258, 245.6, 231.8, 222.8, 216.8, 
    218.6, 214.8, _, _, _, _, _, _, _, _, _, _,
  291.3, -99999, 292.5, 295.7, 284.9, 261.4, 251, 235.4, 225.8, 213.8, 202, 
    206.4, _, _, _, _, _, _, _, _, _, _,
  291.9, -99999, -99999, 298.7, 284.7, 262.2, 251.2, 235.4, 225, 213.6, 
    203.6, 205.6, _, _, _, _, _, _, _, _, _, _,
  288.9, -99999, -99999, -99999, 278.1, 259.6, 250.2, 233.4, 224.6, 212.8, 
    206.2, 210.8, _, _, _, _, _, _, _, _, _, _,
  292.5, -99999, -99999, -99999, 282.3, 260.8, 248.4, 232.8, 223.6, 212.4, 
    212.8, 212.4, _, _, _, _, _, _, _, _, _, _,
  285.1, 283.9, 282.1, 281.5, 271.4, 253.8, 240.2, 227.8, 220.6, 224.2, 
    221.2, 216.4, _, _, _, _, _, _, _, _, _, _,
  291.1, -99999, 292.5, 293.9, 283.7, 261.2, 249.8, 234.8, 224.2, 214.4, 
    205.8, 210.4, _, _, _, _, _, _, _, _, _, _,
  286.9, -99999, -99999, 288.1, 280.9, 261.2, 248.8, 233.8, 224.8, 214, 
    204.4, 210.8, _, _, _, _, _, _, _, _, _, _,
  280.7, -99999, -99999, -99999, 275.1, 253, 241.8, 228.2, 220.2, 219.8, 
    219.8, 216, _, _, _, _, _, _, _, _, _, _,
  290.9, -99999, 289.3, 287.7, 278.5, 262.8, 251.2, 236, 226, 214, 203.8, 
    211.6, _, _, _, _, _, _, _, _, _, _,
  284.7, -99999, 282.1, 280.7, 276.5, 260.6, 247, 233.4, 223.6, 213.6, 210.4, 
    214.2, _, _, _, _, _, _, _, _, _, _,
  282.1, -99999, -99999, 281.7, 271.6, 253.6, 240.4, 225.6, 220.8, 220, 221, 
    216.8, _, _, _, _, _, _, _, _, _, _,
  283.1, -99999, 280.7, 278.1, 270.4, 257.6, 244.8, 231.4, 222.4, 217.6, 
    218.8, 214, _, _, _, _, _, _, _, _, _, _,
  280.5, -99999, 287.1, 283.5, 270.2, 253.4, 241.2, 228.4, 219.2, 216.6, 
    219.2, 218, _, _, _, _, _, _, _, _, _, _,
  280.9, -99999, 282.9, 283.1, 270.4, 254, 241.6, 224.6, 215, 220, 219.6, 
    217.2, _, _, _, _, _, _, _, _, _, _,
  299.9, 300.1, 295.9, 291.5, 283.1, 266.8, 254.4, 239, 229.8, 220, 208.4, 
    197.2, _, _, _, _, _, _, _, _, _, _,
  264, 266.8, 265.8, 262.4, 255.4, 241.8, 230.4, 224, 226.6, 228.8, 230, 
    228.8, _, _, _, _, _, _, _, _, _, _,
  282.5, 281.7, 284.7, 278.3, 269.6, 256, 245.8, 228.4, 218.8, 214, 214.2, 
    215.8, _, _, _, _, _, _, _, _, _, _,
  285.5, -99999, 285.3, 280.7, 274.3, 258.6, 248.8, 232, 222.2, 213.6, 204.6, 
    212.2, _, _, _, _, _, _, _, _, _, _,
  277.7, 275.5, 276.5, 271, 264.8, 250.2, 237.8, 223.6, 218.8, 222.4, 221.4, 
    219, _, _, _, _, _, _, _, _, _, _,
  275.1, 275.1, 274.3, 269.8, 265.4, 249.8, 237, 223, 216, 220.4, 224.8, 
    225.4, _, _, _, _, _, _, _, _, _, _,
  266.4, -99999, 268.2, 270, 265, 249.6, 238, 223.6, 220, 226.8, 225.8, 
    226.6, _, _, _, _, _, _, _, _, _, _,
  291.9, 291.1, 287.3, 284.5, 278.5, 261, 250.6, 233.4, 223.6, 212.2, 204.2, 
    207, _, _, _, _, _, _, _, _, _, _,
  296.9, 296.3, 290.9, 288.3, 280.7, 262.6, 250.4, 235.4, 226.6, 216.6, 
    207.4, 205.8, _, _, _, _, _, _, _, _, _, _,
  290.9, 294.5, 292.1, 286.3, 278.1, 264, 251.4, 234.2, 224, 212.4, 204, 206, 
    _, _, _, _, _, _, _, _, _, _,
  293.1, 294.9, 291.5, 286.9, 277.5, 263, 250.8, 235, 224.6, 213.6, 202.4, 
    208.2, _, _, _, _, _, _, _, _, _, _,
  292.7, 295.1, 292.1, 287.5, 277.1, 262.6, 252, 234.2, 224.6, 213, 202.2, 
    205.2, _, _, _, _, _, _, _, _, _, _,
  287.7, -99999, 292.5, 287.1, 278.3, 263, 251.6, 235.8, 225, 213, 201.6, 
    206.4, _, _, _, _, _, _, _, _, _, _,
  293.7, 295.7, 291.1, 289.7, 280.3, 263.2, -99999, -99999, -99999, -99999, 
    -99999, -99999, _, _, _, _, _, _, _, _, _, _,
  295.9, 294.5, 289.9, 289.5, 283.1, 263.6, 251.8, 236.4, 226, 214.8, 201.6, 
    -99999, _, _, _, _, _, _, _, _, _, _,
  287.3, -99999, 290.7, 287.3, 277.9, 263.6, 252, 233.8, 224.6, 213, 201.2, 
    206.2, _, _, _, _, _, _, _, _, _, _,
  283.7, 286.3, 284.7, 280.7, 274.9, 262.2, 247.8, 230.6, 219.8, 211, 209.4, 
    209.4, _, _, _, _, _, _, _, _, _, _,
  287.1, -99999, 289.3, 284.5, 276.7, 260.8, 250.2, 233.4, 222.6, 211.4, 
    204.4, 210.4, _, _, _, _, _, _, _, _, _, _,
  297.1, 297.7, 292.1, 287.7, 280.7, 265.4, 256.8, 241.6, 232, 219.2, 205.2, 
    199.4, _, _, _, _, _, _, _, _, _, _,
  297.5, 296.9, 292.1, 288.5, 280.1, 266.2, 253.6, 238.4, 229, 218, 207.4, 
    200.8, _, _, _, _, _, _, _, _, _, _,
  296.5, 296.7, 291.9, 288.3, 280.9, 266.4, 254, 237.8, 228.2, 216.2, 207, 
    201.6, _, _, _, _, _, _, _, _, _, _,
  292.1, -99999, -99999, 292.7, 281.7, 261, 251.8, 236.2, 225.8, 213.8, 
    210.8, 207.2, _, _, _, _, _, _, _, _, _, _,
  289.3, -99999, 283.1, 282.5, 277.9, 260.8, 249, 233.6, 224.6, 213.4, 212.4, 
    215, _, _, _, _, _, _, _, _, _, _,
  281.1, -99999, -99999, -99999, 271.2, 252.6, 239.4, 225.4, 222.4, 222.8, 
    222.6, 218.2, _, _, _, _, _, _, _, _, _, _,
  285.9, -99999, -99999, 288.1, 278.9, 257.4, 245, 231.2, 222, 212, 217, 215, 
    _, _, _, _, _, _, _, _, _, _,
  282.5, -99999, 283.7, 280.1, 270.8, 253.4, 240.4, 223, 221, 222.6, 221.2, 
    216.4, _, _, _, _, _, _, _, _, _, _,
  285.5, -99999, 287.7, 287.3, 276.5, 262.2, 250.8, 234.2, 223.6, 212.4, 
    203.8, 211.2, _, _, _, _, _, _, _, _, _, _,
  290.7, -99999, 290.1, 287.9, 277.7, 261.6, 248.8, 233.4, 225, 214, 208.2, 
    212.4, _, _, _, _, _, _, _, _, _, _,
  284.3, -99999, -99999, 281.5, 275.9, 258.2, 246.4, 232.2, 223.4, 213.4, 
    209.2, 213.6, _, _, _, _, _, _, _, _, _, _,
  277.5, -99999, -99999, 282.7, 270.8, 254, 240.6, 226.6, 218.8, 218, 219.4, 
    217.2, _, _, _, _, _, _, _, _, _, _,
  283.1, 283.1, 279.1, 282.1, 272.4, 254.8, 242.4, 227.4, 218, 215.4, 218.6, 
    215.8, _, _, _, _, _, _, _, _, _, _,
  295.1, -99999, 293.9, 290.1, 283.1, 264.2, 251.4, 234.8, 224.2, 213.6, 
    202.6, 211.2, _, _, _, _, _, _, _, _, _, _,
  299.7, 299.5, 294.5, 290.9, 283.3, 268, 257.6, 242.8, 232, 220.8, 206, 
    194.6, _, _, _, _, _, _, _, _, _, _,
  299.9, 299.7, 295.7, 292.5, 282.7, 267.4, 257.4, 242, 232.6, 219.6, 206, 
    193.4, _, _, _, _, _, _, _, _, _, _,
  301.1, 300.7, 296.9, 292.3, 283.3, 267.4, 258.6, 243.4, 233.2, 220.8, 
    206.2, 192, _, _, _, _, _, _, _, _, _, _,
  262.8, 260.8, 268.4, 269.4, 259.2, 243.2, 232.4, 221, 222, 227.8, 228.4, 
    228.6, _, _, _, _, _, _, _, _, _, _,
  280.9, 279.7, 278.3, 273.9, 268.2, 250.8, 240, 227.4, 217.8, 213.8, 217.2, 
    219.4, _, _, _, _, _, _, _, _, _, _,
  279.3, 277.5, 271.8, 266.4, 262.6, 247.6, 234.6, 223.2, 219.2, 223.4, 
    226.2, 225, _, _, _, _, _, _, _, _, _, _,
  271.2, -99999, 267.6, 271.2, 267.8, 253.8, 241.2, 225.8, 218.8, 224.8, 
    219.4, 219.6, _, _, _, _, _, _, _, _, _, _,
  268.2, -99999, 264, 266.6, 260.8, 248.4, 237.4, 222, 219.8, 224.8, 225, 
    220.4, _, _, _, _, _, _, _, _, _, _,
  273.7, 273, 268, 262.8, 260, 245, 232.2, 221.4, 225.6, 228, 228.8, 228.6, 
    _, _, _, _, _, _, _, _, _, _,
  260.4, 264.6, 262, 264.8, 259.4, 242.8, 232.8, 221, 225, 227.8, 227.8, 
    227.6, _, _, _, _, _, _, _, _, _, _,
  267, 267.6, 265.2, 264.2, 259.4, 243.6, 232.2, 219.4, 222.6, 226.2, 226, 
    224.8, _, _, _, _, _, _, _, _, _, _,
  270.8, 269, 271.4, 268, 258.4, 241.8, 230.6, 220.6, 226.4, 228.6, 227.4, 
    224.8, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  275.1, 274.5, 270.8, 268.8, 259.8, 242.2, 231.4, 220, 227.4, 226.4, 228, 
    222.8, _, _, _, _, _, _, _, _, _, _,
  285.3, 286.1, 282.9, 278.3, 268.6, 254.6, 244.4, 227.2, 220.4, 218, 219.8, 
    217.2, _, _, _, _, _, _, _, _, _, _,
  299.7, 299.3, 295.9, -99999, -99999, 267.8, -99999, 243.4, 233.2, 220, 
    203.4, 196.8, _, _, _, _, _, _, _, _, _, _,
  284.1, -99999, 286.1, 282.7, 272.6, 253.4, 240.6, 225, 216, 220, 219.4, 
    217.6, _, _, _, _, _, _, _, _, _, _,
  280.3, 282.7, 279.7, 274.3, 271, 255.2, 243.4, 228.8, 219.8, 215.4, 215.4, 
    216, _, _, _, _, _, _, _, _, _, _,
  265.6, 264.4, 271.6, 269.4, 261.8, 245, 233.4, 221.2, 221.4, 229, 226.4, 
    227.8, _, _, _, _, _, _, _, _, _, _,
  260, 258.4, 254.4, 262, 258.8, 243.2, 232.4, 219.2, 222, 228.2, 230.2, 
    228.2, _, _, _, _, _, _, _, _, _, _,
  297.5, 297.3, 292.5, 287.9, 285.5, 268.6, 254.6, 241.2, 231.6, 219.8, 
    207.6, 196.6, _, _, _, _, _, _, _, _, _, _,
  282.5, 281.7, 283.7, 285.1, 273, 256.8, 244, 227.8, 219.6, 210.2, 217.2, 
    214.8, _, _, _, _, _, _, _, _, _, _,
  279.9, -99999, 279.5, 274.7, 266.4, 251, 237.6, 222, 213.8, 221.6, 222.2, 
    218.4, _, _, _, _, _, _, _, _, _, _,
  297.5, 297.3, 293.9, 288.7, 282.9, 266.8, 255.4, 243.4, 233.4, 219.6, 
    205.2, 196.4, _, _, _, _, _, _, _, _, _, _,
  296.1, -99999, 294.3, 291.1, 279.5, 261.4, 249.4, 234.4, 225, 213.8, 
    -99999, -99999, _, _, _, _, _, _, _, _, _, _,
  297.9, 297.5, -99999, 289.9, 281.1, -99999, -99999, -99999, -99999, 219.2, 
    204.4, 199.8, _, _, _, _, _, _, _, _, _, _,
  278.7, 276.7, 276.9, 273.7, 265.2, 250, 238.2, 222.8, 214.8, 222.6, -99999, 
    -99999, _, _, _, _, _, _, _, _, _, _,
  285.1, 285.3, 280.9, 284.5, 275.3, 258, 246.4, 232.6, 224, 218, -99999, 
    -99999, _, _, _, _, _, _, _, _, _, _,
  285.3, -99999, -99999, 283.5, 276.1, 257, 245.8, 229.6, 225, 219.2, 218, 
    216.6, _, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 0, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 0, _, _, _, _, _, _, _, _, _,
  296.5, 296.9, 293.7, 289.9, 281.3, 268, 258, 240.8, 230.8, 218.8, 205.6, 
    194.6, _, _, _, _, _, _, _, _, _, _ ;

 tdMan =
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 1.249117e-40, _, _, _, _, _, _, _, _, _,
  2.600006, -99999, -99999, 4.200012, 17, 18.99998, 15, 12, -99999, -99999, 
    -99999, -99999, _, _, _, _, _, _, _, _, _, _,
  1.200012, 3.399994, 2.299988, 1.700012, 2.300003, 3.600006, 5, 8, 16, 29, 
    29, 28, _, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 1.249117e-40, _, _, _, _, _, _, _, _, _,
  2.100006, -99999, 0.6000061, 15, 38, 32, 29, 23, 22, 22, 21, 20, 
    1.249117e-40, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 1.249117e-40, _, _, _, _, _, _, _, _, _,
  0.7000122, 2, 2.299988, 2.200012, 3.399994, 11, 12, 5, 5, 4.199997, 7, 6, 
    _, _, _, _, _, _, _, _, _, _,
  1.5, -99999, 2.600006, 0.6999817, 1.199982, 10, 10, 7, 10, 34, 34, 33, _, 
    _, _, _, _, _, _, _, _, _,
  0, 0.2999878, 6, 4.800018, 3.5, 10, 11, 9, 11, 21, 23, 24, _, _, _, _, _, 
    _, _, _, _, _,
  0, 0.7000122, 0.8999939, 1, 1, 2.400009, 3.699997, 5, 6, 6, 8, 12, _, _, _, 
    _, _, _, _, _, _, _,
  1.200012, 1.700012, 1.900024, 3, 0.3000183, 2.300003, 3, 3.199997, 
    3.399994, 3.099991, 6, 15, _, _, _, _, _, _, _, _, _, _,
  1.5, 2.700012, 0.7999878, 13, 19, 4.300003, 3.900009, 3.699997, 4, 
    4.100006, 8, 23, _, _, _, _, _, _, _, _, _, _,
  1.700012, 2.899994, 12, 18, 21, 4.100006, 3.100006, 7, 4.600006, 4.800003, 
    7, 20, _, _, _, _, _, _, _, _, _, _,
  3.200012, 2.5, 2, 2.899994, 12, 7, 15, 6, 17, 13, 12, 11, _, _, _, _, _, _, 
    _, _, _, _,
  1.399994, 3.200012, 3.799988, 4.299988, 6, 6, 6.000015, 3.200012, 4.5, 5, 
    4.899994, 5, _, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 1.249117e-40, _, _, _, _, _, _, _, _, _,
  1.800018, 1.399994, 2.300018, 0.9000244, 4, 8, 11, 9, 18, 23, 24, 23, _, _, 
    _, _, _, _, _, _, _, _,
  2.800018, 11, 5, 0.7000122, 12, 1.699997, 4.5, 6, 5, 3.5, 14, 25, _, _, _, 
    _, _, _, _, _, _, _,
  1.700012, 7, 7, 2.100006, 8, 13, 7, 7, 6, 4.400009, 20, 23, _, _, _, _, _, 
    _, _, _, _, _,
  4.399994, 7, 10, 3.799988, 0.6000061, 10, 10, 10, 12, 18, 23, 23, _, _, _, 
    _, _, _, _, _, _, _,
  2.200012, 5, 4.899994, 4, 6, 2.799988, 4.900009, 2.800003, 3, 3.699997, 15, 
    22, _, _, _, _, _, _, _, _, _, _,
  0, 0.6999817, 4.399994, 18, 14, 4.600006, 4.599991, 3.5, 3.300003, 
    3.199997, 16, 23, _, _, _, _, _, _, _, _, _, _,
  3.300018, 5, 9, 8, 19, 7, 8, 5, 5, 5, 6, 8, _, _, _, _, _, _, _, _, _, _,
  1.699982, 3.800018, 0.7999878, 3, 4.899994, 7, 10, 3.199997, 9, 8, 10, 9, 
    _, _, _, _, _, _, _, _, _, _,
  2.900024, 3.099976, 2.400024, 1.5, 6, 3.399994, 1.5, 4.199997, 10, 8, 
    4.399994, 4.100006, _, _, _, _, _, _, _, _, _, _,
  1.5, 3.699982, 7, 4.700012, 28, 23, 28, 19, 10, 8, 8, 12, _, _, _, _, _, _, 
    _, _, _, _,
  2.699982, -99999, -99999, -99999, 1, 2.5, 6, 3.699997, 2.899994, 4, 12, 19, 
    _, _, _, _, _, _, _, _, _, _,
  2.200012, -99999, 1.100006, 0.8999939, 25.99998, 16, 9, 9, 8, 8, 9, 13, _, 
    _, _, _, _, _, _, _, _, _,
  0.9000244, 2.700012, 4.600006, 4.299988, 6, 6, 5, 18, 2.699997, 3.100006, 
    4.399994, 5, _, _, _, _, _, _, _, _, _, _,
  3, 4.099976, 7, 6, 29, 27, 22, 14, 14, 20, 29, 33, _, _, _, _, _, _, _, _, 
    _, _,
  1.199982, 2, 3.600006, 0.6000061, 4.700012, 6, 4.199997, 8, 26, 36, 36, 36, 
    _, _, _, _, _, _, _, _, _, _,
  3.799988, 4.700012, 3.900024, 7, 34.00002, 23.00002, 17, 19, 17, 12, 12, 
    15, _, _, _, _, _, _, _, _, _, _,
  1.199982, 0.5999756, 6, 11, 11, 24, 21, 19, 14, 11, 9, 10, _, _, _, _, _, 
    _, _, _, _, _,
  2.100006, 3, 5, 3.599976, 6, 7, 24, 17, 10, 6, 4.899994, 12, _, _, _, _, _, 
    _, _, _, _, _,
  0, -99999, 6, 5, 4.799988, 12.00002, 25, 14, 7, 7, 5, 11, _, _, _, _, _, _, 
    _, _, _, _,
  1.200012, 1.200012, 2.100006, 3.899994, 5, 7, 12, 8, 4.299988, 7, 6, 7, _, 
    _, _, _, _, _, _, _, _, _,
  0.8000183, 0.5, 1, 3.800018, 8, 42, 37, 5, 6, 5, 4.899994, 12, _, _, _, _, 
    _, _, _, _, _, _,
  0.3000183, -99999, 1.700012, 1.600006, 3.599976, 12, 9, 9, 8, 4.699997, 
    4.5, 9, _, _, _, _, _, _, _, _, _, _,
  1.699982, 0.8999939, 8, 8, 14, 11, 4.600006, 4.800003, 3.900009, 3.600006, 
    3.700012, 23, _, _, _, _, _, _, _, _, _, _,
  0.3000183, -99999, 2.800018, 3, 1.600006, 37.00002, 13, 13, 9, 8, 7, 8, _, 
    _, _, _, _, _, _, _, _, _,
  3.599976, -99999, 0.7999878, 0.5, 13, 1.299988, 2.100006, 2.900009, 3.5, 
    3.300003, 4.100006, 7, _, _, _, _, _, _, _, _, _, _,
  2.400024, 2.5, 14, 11, 18.00002, 16, 4.5, 5, 6, 6, 7, 8, _, _, _, _, _, _, 
    _, _, _, _,
  5, 11, 14, 9, 21, 31.00002, 11, 10, 9, 6, 11, 19, _, _, _, _, _, _, _, _, 
    _, _,
  3.299988, 14, 14, 13, 31.00002, 28.99998, 16, 16, 11, 7, 11, 17, _, _, _, 
    _, _, _, _, _, _, _,
  1.399994, -99999, 3.200012, 1.200012, 25, 28, 19, 16, 8, 6, 4.699997, 10, 
    _, _, _, _, _, _, _, _, _, _,
  1.199982, 1.200012, 6, 14, 7, 7.000015, 16, 19, 16, 12, 9, 15, _, _, _, _, 
    _, _, _, _, _, _,
  2.399994, -99999, 5, 9, 23, 33, 30, 14, 13, 11, 8, 12, _, _, _, _, _, _, _, 
    _, _, _,
  2.299988, -99999, 0.7000122, 0.7000122, -99999, -99999, -99999, 29, 18, 13, 
    11, 10, _, _, _, _, _, _, _, _, _, _,
  2.799988, -99999, -99999, 1.299988, 31, 31.00002, 29, 22, 13, 8, 10, 13, _, 
    _, _, _, _, _, _, _, _, _,
  0.7000122, -99999, 6, 5, 12, 8, 15, -99999, -99999, -99999, -99999, -99999, 
    _, _, _, _, _, _, _, _, _, _,
  2.199982, -99999, 4.299988, 26, 22, 27.99998, 26, 8, 16, 10, 6, 11, _, _, 
    _, _, _, _, _, _, _, _,
  3.800018, -99999, -99999, 6, 21, 16, 19, 14, 8, 6, 5, 11, _, _, _, _, _, _, 
    _, _, _, _,
  14, -99999, -99999, 16, 21, 15, 33, 12, 12, 12, 11, 14, _, _, _, _, _, _, 
    _, _, _, _,
  24, -99999, -99999, -99999, 19, 3.399994, 13, 9, 8, 7, 7, 7, _, _, _, _, _, 
    _, _, _, _, _,
  6, -99999, -99999, -99999, 10, 6, 10, 1.300003, 2.599991, 2.700012, 4, 14, 
    _, _, _, _, _, _, _, _, _, _,
  20, -99999, -99999, 19, 20.99998, 19, 12, 10, 9, 8, 9, 9, _, _, _, _, _, _, 
    _, _, _, _,
  0.5, -99999, 2.200012, 26, 14, 21, 28, 9, 10, 5, 6, 11, _, _, _, _, _, _, 
    _, _, _, _,
  6, -99999, -99999, 19, 13, 2.700012, 15, 4.799988, 5, 6, 5, 6, _, _, _, _, 
    _, _, _, _, _, _,
  10, -99999, -99999, -99999, 3.600006, 3.700012, 24, 3.099991, 2.600006, 
    3.800003, 4.399994, 14, _, _, _, _, _, _, _, _, _, _,
  25, -99999, -99999, -99999, 13, 5.999985, 3.699997, 7, 6, 7, 11, 18, _, _, 
    _, _, _, _, _, _, _, _,
  2.600006, 1.699982, 3.200012, 9, 42, 37, 33, 25, 20, 27, 27, 25, _, _, _, 
    _, _, _, _, _, _, _,
  0.2000122, -99999, 2, 14, 13, 3.300018, 15, 4.900009, 5, 7, 7, 14, _, _, _, 
    _, _, _, _, _, _, _,
  7, -99999, -99999, 14, 11, 7.000015, 22, 12, 15, 4.300003, 4.399994, 15, _, 
    _, _, _, _, _, _, _, _, _,
  6, -99999, -99999, -99999, 8, 3, 13, 11, 10, 10, 10, 10, _, _, _, _, _, _, 
    _, _, _, _,
  0.6999817, -99999, 1, 1.600006, 9, 16.99998, 29, 20, 16, 11, 9, 12, _, _, 
    _, _, _, _, _, _, _, _,
  2.800018, -99999, 2.399994, 3.600006, 15, 18, 1.800003, 13, 11, 8, 10, 19, 
    _, _, _, _, _, _, _, _, _, _,
  3.100006, -99999, -99999, 8, 11, 31, 17, 23, 27, -99999, -99999, -99999, _, 
    _, _, _, _, _, _, _, _, _,
  1.100006, -99999, 1.200012, 2.700012, 8, 28, 16, 16, 10, 14, 22, 22, _, _, 
    _, _, _, _, _, _, _, _,
  0.8999939, -99999, 7, 11, 8, 11, 2.599991, 12, 9, 9, 11, 12, _, _, _, _, _, 
    _, _, _, _, _,
  1.399994, -99999, 2.699982, 8, 1.399994, 6, 12, 12, 9, 13, 24, 25, _, _, _, 
    _, _, _, _, _, _, _,
  2.299988, 2, 3.100006, 3.700012, 8, 9, 8, 9, 11, 11, 9, 7, _, _, _, _, _, 
    _, _, _, _, _,
  1.799988, 0.7999878, 2.699982, 3.299988, 3.799988, 7, 7, 14, 22, 31, 31, 
    31, _, _, _, _, _, _, _, _, _, _,
  1.899994, 2.200012, 15, 9, 16, 23, 29, 11, 10, 10, 18, 25, _, _, _, _, _, 
    _, _, _, _, _,
  5, -99999, 12, 12, 24.99998, 1.800018, 8, 6, 6, 6, 8, 19, _, _, _, _, _, _, 
    _, _, _, _,
  1.800018, 0.1000061, 9, 9, 21.99998, 23, 16, 10, 11, 22, 29, 28, _, _, _, 
    _, _, _, _, _, _, _,
  8, 7, 8, 4.699982, 1.799988, 3.199997, 4, 5, 4, 17, 27, 27, _, _, _, _, _, 
    _, _, _, _, _,
  1.399994, -99999, 0, 27, 2.399994, 2.5, 2.600006, 6, 7, 17, 18, 22, _, _, 
    _, _, _, _, _, _, _, _,
  1.199982, 1.100006, 0, 0, 7, 11, 10, 7, 6, 6, 5, 10, _, _, _, _, _, _, _, 
    _, _, _,
  3.199982, 3.599976, 2.299988, 12, 29.00002, 10, 10, 11, 11, 10, 8, 8, _, _, 
    _, _, _, _, _, _, _, _,
  0.6999817, 2.399994, 13, 1.299988, 7, 23, 20, 10, 9, 7, 6, 12, _, _, _, _, 
    _, _, _, _, _, _,
  0, 0.6999817, 3.899994, 1.600006, 2.100006, 8, 10, 12, 16, 13, 11, 18, _, 
    _, _, _, _, _, _, _, _, _,
  0.8000183, 3, 4.800018, 5, 2.5, 5, 10, 13, 11, 10, 7, 12, _, _, _, _, _, _, 
    _, _, _, _,
  0, -99999, 3.799988, 2.600006, 4.199982, 18, 23, 8, 12, 8, 8, 13, _, _, _, 
    _, _, _, _, _, _, _,
  0.7000122, 2.600006, 3.700012, 11, 19, 15.00002, -99999, -99999, -99999, 
    -99999, -99999, -99999, _, _, _, _, _, _, _, _, _, _,
  1.699982, 1.200012, 0, 9, 23, 32, 17, 18, 13, 9, 7, -99999, _, _, _, _, _, 
    _, _, _, _, _,
  0.5, -99999, 3.5, 2.5, 4.399994, 21, 17, 4.100006, 11, 6, 4.599991, 10, _, 
    _, _, _, _, _, _, _, _, _,
  0.6000061, 4.899994, 13, 22, 36, 22.00002, 22, 4.300003, 3.300003, 
    4.199997, 9, 17, _, _, _, _, _, _, _, _, _, _,
  3.600006, -99999, 3.699982, 7, 29.00002, 12.99998, 8, 3.899994, 3.700012, 
    4.899994, 7, 15, _, _, _, _, _, _, _, _, _, _,
  1.600006, 2.200012, 0.8000183, 0.8000183, 6, 1.100006, 12.99998, 16, 11, 8, 
    7, 7, _, _, _, _, _, _, _, _, _, _,
  2.100006, 1.399994, 1.5, 9, 16, 34.00002, 28, 22, 18, 14, 11, 10, _, _, _, 
    _, _, _, _, _, _, _,
  1.700012, 1.400024, 1.5, 6, 32, 33, 28, 21, 18, 13, 11, 10, _, _, _, _, _, 
    _, _, _, _, _,
  17, -99999, -99999, 21, 21, 16, 28, 12, 6, 6, 11, 16, _, _, _, _, _, _, _, 
    _, _, _,
  5, -99999, 0.7000122, 46, 24, 38.99998, 17, 20, 17, 13, 13, 16, _, _, _, _, 
    _, _, _, _, _, _,
  7, -99999, -99999, -99999, 2.600006, 21, 13, 11, 17, 23, 26, 24, _, _, _, 
    _, _, _, _, _, _, _,
  10, -99999, -99999, 13, 18, 3.299988, 3.300003, 8, 11, 7, 17, 22, _, _, _, 
    _, _, _, _, _, _, _,
  1.600006, -99999, 6, 1.399994, 5, 3.5, 4.599991, 5, 8, 17, 27, 25, _, _, _, 
    _, _, _, _, _, _, _,
  0.6000061, -99999, 0, 4.699982, 1.200012, 5, 13, 2.899994, 3.400009, 3.5, 
    3.699997, 12, _, _, _, _, _, _, _, _, _, _,
  1.200012, -99999, 6, 14, 20, 9, 9, 13, 5, 6, 6, 18, _, _, _, _, _, _, _, _, 
    _, _,
  6, -99999, -99999, 4.299988, 11, 1, 2.699997, 5, 8, 8, 9, 18, _, _, _, _, 
    _, _, _, _, _, _,
  1.100006, -99999, -99999, 7, 2, 11, 7, 11, 11, 11, 16, 20, _, _, _, _, _, 
    _, _, _, _, _,
  1.100006, 1.700012, 1, 5, 13, 20, 33, 9, 8, 8, 11, 12, _, _, _, _, _, _, _, 
    _, _, _,
  1, -99999, 2.399994, 1.200012, 17, 28.00002, 29, 17, 10, 7, 4.900009, 13, 
    _, _, _, _, _, _, _, _, _, _,
  2.300018, 2.100006, 0.5, 0.5, 3.5, 4.5, 38, 33, 6, 8, 7, 6, _, _, _, _, _, 
    _, _, _, _, _,
  2.5, 3.100006, 4.900024, 11, 6, 10, 10, 7, 14, 8, 8, 4.899994, _, _, _, _, 
    _, _, _, _, _, _,
  2.700012, 2.600006, 1.5, 1.399994, 2.899994, 30, 30, 30, 30, -99999, 
    -99999, -99999, _, _, _, _, _, _, _, _, _, _,
  0.8999939, 0, 11, 23, 5.000015, 12, 7, 4.600006, 8, 24, 35, 36, _, _, _, _, 
    _, _, _, _, _, _,
  8, 7, 10, 10, 4.100006, 6, 5, 6, 6, 7, 21, 29, _, _, _, _, _, _, _, _, _, _,
  7, 9, 7, 3.399994, 12, 11, 4.200012, 10, 9, 25, 35, 34, _, _, _, _, _, _, 
    _, _, _, _,
  1.400024, -99999, 0.3000183, 0, 14.99998, 15, 14, 12, 11, 24, 26, 26, _, _, 
    _, _, _, _, _, _, _, _,
  5, -99999, 5, 14, 16.99998, 10, 13, 7, 10, 17, 23, 24, _, _, _, _, _, _, _, 
    _, _, _,
  3.400024, 4.299988, 3.200012, 0.2999878, 10, 18, 8, 10, 22, 31, 31, 31, _, 
    _, _, _, _, _, _, _, _, _,
  3.799988, 2.5, 0.5, 7, 7, 16, 12, 9, 20, 28, 31, 31, _, _, _, _, _, _, _, 
    _, _, _,
  3.899994, 6, 7, 12.00002, 16, 8, 12, 5, 13, 24, 28, 27, _, _, _, _, _, _, 
    _, _, _, _,
  0, 0, 1.899994, 4.600006, 8, 6, 2.5, 4.5, 16, 19, 19, 18, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.200012, 1.600006, 0.6999817, 1.5, 2.099976, 9, 7, 5, 23, 30, 35, 34, _, 
    _, _, _, _, _, _, _, _, _,
  6, 8, 7, 4.799988, 0.7000122, 3.800003, 3.599991, 2.5, 6, 10, 11, 9, _, _, 
    _, _, _, _, _, _, _, _,
  2.700012, 2.699982, 3.399994, -99999, -99999, 11, -99999, 4.699997, 6, 
    -99999, -99999, -99999, _, _, _, _, _, _, _, _, _, _,
  3.100006, -99999, 7, 6, 4.399994, 16, 7, 4, 2.699997, 12, 21, 24, _, _, _, 
    _, _, _, _, _, _, _,
  4.699982, 9, 16, 13, 28, 22, 23, 20, 5, 11, 19, 28, _, _, _, _, _, _, _, _, 
    _, _,
  3, 4.799988, 14, 17, 21.99998, 16, 12, 11, 15, 36, 35, 35, _, _, _, _, _, 
    _, _, _, _, _,
  2, 3.099991, 0.1999969, 6, 15.99998, 8, 10, 6, 10, 19, 27, 28, _, _, _, _, 
    _, _, _, _, _, _,
  3.299988, 4.899994, 5, 9, 27, 26, 3.600006, 13, -99999, -99999, -99999, 
    -99999, _, _, _, _, _, _, _, _, _, _,
  2.100006, 0.8000183, 8, 19, 20, 8.999985, 8, 5, 4.400009, 4.099991, 17, 31, 
    _, _, _, _, _, _, _, _, _, _,
  7, -99999, 8, 5, 2.299988, 7, 2.900009, 3.800003, 4, 23, 27, 26, _, _, _, 
    _, _, _, _, _, _, _,
  1, 1.099976, 1.100006, 1.200012, 3.399994, 0.8999939, 8, 7, 9, 11, 11, 9, 
    _, _, _, _, _, _, _, _, _, _,
  26, -99999, 29, 22, 16, 13, 9, 7, -99999, -99999, -99999, -99999, _, _, _, 
    _, _, _, _, _, _, _,
  6, 6, -99999, 6, 8, -99999, -99999, -99999, -99999, 8, 7, 7, _, _, _, _, _, 
    _, _, _, _, _,
  2.800018, 2.800018, 8, 3.600006, 2.400024, 7, 10, -99999, -99999, -99999, 
    -99999, -99999, _, _, _, _, _, _, _, _, _, _,
  4.300018, 3.5, 2.699982, 11, 28.99998, 40, 24, -99999, -99999, -99999, 
    -99999, -99999, _, _, _, _, _, _, _, _, _, _,
  7, -99999, -99999, 11, 33, 29, 26, 20, 19, 17, 17, 17, _, _, _, _, _, _, _, 
    _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 1.249117e-40, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 1.249117e-40, _, _, _, _, _, _, _, _, _,
  1.600006, 1.699982, 3, 4.699982, 3.199982, 34, 33, 28, -99999, -99999, 
    -99999, -99999, _, _, _, _, _, _, _, _, _, _ ;

 wdMan =
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 0, _, _, _, _, _, _, _, _, _,
  50, 60, -99999, 85, 90, 70, 310, 5, 265, 265, 250, 270, _, _, _, _, _, _, 
    _, _, _, _,
  180, 190, 210, 225, 225, 245, 245, 250, 255, 245, 245, 300, _, _, _, _, _, 
    _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 0, _, _, _, _, _, _, _, _, _,
  325, -99999, 345, 10, 270, 260, 255, 245, 235, 240, 255, 230, 0, _, _, _, 
    _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 0, _, _, _, _, _, _, _, _, _,
  130, 120, 225, 215, 80, 55, 65, 105, 125, 190, 225, 250, _, _, _, _, _, _, 
    _, _, _, _,
  60, -99999, 100, 200, 335, 295, 305, 310, 320, 325, 325, 330, _, _, _, _, 
    _, _, _, _, _, _,
  90, 155, 200, 205, 245, 245, 245, 245, 245, 240, 240, 225, _, _, _, _, _, 
    _, _, _, _, _,
  80, -99999, -99999, 130, 115, 175, 175, 190, 195, 190, 200, 190, _, _, _, 
    _, _, _, _, _, _, _,
  140, 140, 145, 165, 180, 170, 185, 180, 175, 180, 180, 195, _, _, _, _, _, 
    _, _, _, _, _,
  250, 260, 85, 160, 215, 240, 245, 250, 250, 265, 255, 255, _, _, _, _, _, 
    _, _, _, _, _,
  320, 315, 230, 250, 245, 255, 245, 260, 275, 280, 270, 275, _, _, _, _, _, 
    _, _, _, _, _,
  190, 190, 195, 195, 245, 260, 280, 250, 260, 265, 265, 260, _, _, _, _, _, 
    _, _, _, _, _,
  170, 165, 155, 160, 155, 140, 50, 320, 340, 15, 30, 355, _, _, _, _, _, _, 
    _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 0, _, _, _, _, _, _, _, _, _,
  230, 240, 240, 245, 240, 240, 250, 250, 245, 240, 240, 230, _, _, _, _, _, 
    _, _, _, _, _,
  340, 30, 125, 205, 245, 240, 245, 245, 240, 245, 240, 240, _, _, _, _, _, 
    _, _, _, _, _,
  300, 320, 45, 255, 260, 265, 265, 265, 265, 265, 260, 250, _, _, _, _, _, 
    _, _, _, _, _,
  40, 25, 235, 255, 270, 275, 275, 285, 285, 280, 285, 295, _, _, _, _, _, _, 
    _, _, _, _,
  150, 225, 340, 5, 280, 270, 275, 270, 280, 280, 275, 280, _, _, _, _, _, _, 
    _, _, _, _,
  140, 145, 320, 320, 295, 305, 305, 305, 300, 305, 310, 320, _, _, _, _, _, 
    _, _, _, _, _,
  340, 345, 10, 355, 325, 330, 325, 330, 335, 325, 330, 345, _, _, _, _, _, 
    _, _, _, _, _,
  200, -99999, 320, 190, 245, 275, 285, 255, 240, 235, 275, 230, _, _, _, _, 
    _, _, _, _, _, _,
  30, 30, 360, 335, 90, 75, 110, 120, 140, 200, 205, 250, _, _, _, _, _, _, 
    _, _, _, _,
  100, 115, 105, 60, 35, 65, 50, 50, 40, 15, 335, 310, _, _, _, _, _, _, _, 
    _, _, _,
  85, -99999, -99999, -99999, 155, 235, 215, 225, 220, 225, 230, 235, _, _, 
    _, _, _, _, _, _, _, _,
  350, -99999, 40, 10, 335, 275, 260, 255, 255, 250, 250, 265, _, _, _, _, _, 
    _, _, _, _, _,
  120, 105, 65, 45, 60, 360, 315, 245, 220, 225, 260, 300, _, _, _, _, _, _, 
    _, _, _, _,
  330, 340, 360, 360, 290, 255, 245, 250, 250, 245, 255, 220, _, _, _, _, _, 
    _, _, _, _, _,
  355, 5, 5, 5, 5, 20, 60, 40, 20, 15, 360, 45, _, _, _, _, _, _, _, _, _, _,
  90, 90, 90, 70, 70, 40, 20, 40, 20, 275, 280, 295, _, _, _, _, _, _, _, _, 
    _, _,
  0, 315, 205, 200, 110, 20, 35, 35, 45, 45, 30, 305, _, _, _, _, _, _, _, _, 
    _, _,
  240, 250, 285, 285, 305, 325, 30, 355, 360, 5, 360, 310, _, _, _, _, _, _, 
    _, _, _, _,
  0, -99999, 305, 300, 290, 300, 350, 320, 345, 5, 355, 310, _, _, _, _, _, 
    _, _, _, _, _,
  185, 185, 250, 275, 300, 340, 15, 295, 275, 320, 345, 300, _, _, _, _, _, 
    _, _, _, _, _,
  60, 75, 75, 315, 295, 315, 290, 315, 335, 350, 340, 315, _, _, _, _, _, _, 
    _, _, _, _,
  210, -99999, 255, 245, 270, 300, 285, 300, 295, 305, 320, 285, _, _, _, _, 
    _, _, _, _, _, _,
  175, 175, 175, 150, 235, 290, 300, 300, 320, 340, 320, 300, _, _, _, _, _, 
    _, _, _, _, _,
  155, -99999, 215, 250, 255, 285, 285, 300, 310, 325, 315, 300, _, _, _, _, 
    _, _, _, _, _, _,
  230, -99999, 245, 260, 250, 260, 280, 280, 290, 290, 300, 285, _, _, _, _, 
    _, _, _, _, _, _,
  0, -99999, 225, 295, 295, 310, 310, 315, 325, 325, 305, 285, _, _, _, _, _, 
    _, _, _, _, _,
  340, 25, 145, 180, 305, 330, 310, 315, 325, 330, 315, 300, _, _, _, _, _, 
    _, _, _, _, _,
  350, 30, 85, 70, 345, 330, 330, 325, 330, 330, 315, 310, _, _, _, _, _, _, 
    _, _, _, _,
  190, -99999, 260, 265, 270, 275, 285, 285, 285, 275, 280, 270, _, _, _, _, 
    _, _, _, _, _, _,
  120, 170, 190, 160, 70, 50, 80, 55, 60, 45, 40, 320, _, _, _, _, _, _, _, 
    _, _, _,
  170, -99999, 200, 195, 130, 45, 235, 235, 265, 225, 290, 295, _, _, _, _, 
    _, _, _, _, _, _,
  135, -99999, -99999, 165, 240, 240, 170, 275, 280, 295, 280, 290, _, _, _, 
    _, _, _, _, _, _, _,
  150, -99999, -99999, 180, 145, 190, 220, 245, 240, 260, 265, 280, _, _, _, 
    _, _, _, _, _, _, _,
  210, -99999, 235, 230, 170, 35, 30, 265, -99999, -99999, 250, 310, _, _, _, 
    _, _, _, _, _, _, _,
  190, -99999, 210, 220, 170, 270, 245, 225, 230, 230, 265, 285, _, _, _, _, 
    _, _, _, _, _, _,
  235, -99999, -99999, 220, 180, 195, 205, 220, 230, 225, 255, 290, _, _, _, 
    _, _, _, _, _, _, _,
  150, -99999, -99999, 175, 275, 230, 230, 235, 235, 250, 240, 240, _, _, _, 
    _, _, _, _, _, _, _,
  220, -99999, -99999, -99999, 225, 220, 225, 225, 230, 235, 245, 250, _, _, 
    _, _, _, _, _, _, _, _,
  220, -99999, -99999, -99999, 215, 215, 215, 215, 225, 225, 230, 220, _, _, 
    _, _, _, _, _, _, _, _,
  190, -99999, -99999, 195, 185, 210, 210, 210, 215, 220, 220, 210, _, _, _, 
    _, _, _, _, _, _, _,
  180, -99999, 230, 255, 290, 300, 240, 280, 285, 275, 240, 285, _, _, _, _, 
    _, _, _, _, _, _,
  190, -99999, -99999, 225, 255, 215, 235, 230, 220, 240, 250, 260, _, _, _, 
    _, _, _, _, _, _, _,
  10, -99999, -99999, -99999, 110, 220, 235, 225, 220, 220, 240, 265, _, _, 
    _, _, _, _, _, _, _, _,
  130, -99999, -99999, -99999, 235, 205, 225, 225, 225, 225, 225, 265, _, _, 
    _, _, _, _, _, _, _, _,
  210, 215, 285, 305, 280, 250, 235, 260, 255, 245, 255, 260, _, _, _, _, _, 
    _, _, _, _, _,
  340, -99999, -99999, 10, 255, 255, 240, 245, 245, 255, 250, 255, _, _, _, 
    _, _, _, _, _, _, _,
  360, -99999, -99999, 30, 160, 235, 245, 240, 240, 240, 240, 250, _, _, _, 
    _, _, _, _, _, _, _,
  130, -99999, -99999, -99999, 70, 200, 200, 205, 210, 215, 215, 230, _, _, 
    _, _, _, _, _, _, _, _,
  240, -99999, 275, 285, 290, 280, 280, 260, 255, 255, 275, 275, _, _, _, _, 
    _, _, _, _, _, _,
  360, -99999, 15, 345, 325, 270, 255, 260, 255, 255, 255, 260, _, _, _, _, 
    _, _, _, _, _, _,
  100, -99999, -99999, 295, 205, 215, 215, 215, 215, 215, 225, 235, _, _, _, 
    _, _, _, _, _, _, _,
  330, -99999, 355, 355, 340, 280, 265, 265, 270, 260, 270, 265, _, _, _, _, 
    _, _, _, _, _, _,
  90, -99999, 100, 115, 320, 275, 260, 250, 245, 250, 245, 260, _, _, _, _, 
    _, _, _, _, _, _,
  10, -99999, 15, 70, 55, 70, 10, 30, 55, 280, 265, 270, _, _, _, _, _, _, _, 
    _, _, _,
  80, 80, 100, 65, 5, 315, 5, 300, 280, 335, 5, 35, _, _, _, _, _, _, _, _, 
    _, _,
  360, 65, 80, 85, 85, 85, 65, 80, 90, 95, 90, 85, _, _, _, _, _, _, _, _, _, _,
  0, 185, 60, 35, 340, 335, 330, 340, 350, 330, 305, 305, _, _, _, _, _, _, 
    _, _, _, _,
  160, -99999, 195, 190, 225, 260, 275, 295, 300, 305, 290, 295, _, _, _, _, 
    _, _, _, _, _, _,
  210, 245, 325, 330, 325, 320, 315, 315, 285, 290, 270, 255, _, _, _, _, _, 
    _, _, _, _, _,
  150, 150, 180, 205, 240, 280, 275, 280, 290, 280, 285, 295, _, _, _, _, _, 
    _, _, _, _, _,
  295, -99999, 280, 250, 230, 230, 225, 235, 235, 255, 255, 255, _, _, _, _, 
    _, _, _, _, _, _,
  90, 100, 130, 260, 290, 290, 305, 320, 345, 355, 330, 305, _, _, _, _, _, 
    _, _, _, _, _,
  60, 75, 90, 75, 80, 340, 310, 340, 280, 270, 265, 285, _, _, _, _, _, _, _, 
    _, _, _,
  210, 190, 190, 35, 65, 345, 345, 25, 30, 20, 20, 320, _, _, _, _, _, _, _, 
    _, _, _,
  210, 220, 250, 325, 90, 315, 330, 20, 35, 40, 25, 285, _, _, _, _, _, _, _, 
    _, _, _,
  0, 115, 20, -99999, -99999, 40, 70, 360, 40, 45, 15, 330, _, _, _, _, _, _, 
    _, _, _, _,
  270, -99999, 295, 300, 15, 355, 40, 30, 30, 30, 45, 335, _, _, _, _, _, _, 
    _, _, _, _,
  190, 185, 175, 170, 145, 75, -99999, -99999, -99999, -99999, -99999, 
    -99999, _, _, _, _, _, _, _, _, _, _,
  180, 190, 210, 195, 120, 110, 35, 360, 20, 290, 245, -99999, _, _, _, _, _, 
    _, _, _, _, _,
  0, -99999, 285, 305, 285, 320, 330, 305, 350, 10, 350, 310, _, _, _, _, _, 
    _, _, _, _, _,
  360, 35, 105, 95, 305, 305, 300, 305, 310, 330, 325, 310, _, _, _, _, _, _, 
    _, _, _, _,
  160, -99999, -99999, 240, 250, 270, 285, 310, 305, 315, 305, 295, _, _, _, 
    _, _, _, _, _, _, _,
  130, 110, 95, 90, 135, 250, 255, 275, 255, 255, 275, 285, _, _, _, _, _, _, 
    _, _, _, _,
  140, 145, 160, 150, 120, 20, 15, 305, 305, 305, 305, 310, _, _, _, _, _, _, 
    _, _, _, _,
  140, 145, 160, 160, 140, 40, 15, 310, 305, 305, 310, 315, _, _, _, _, _, _, 
    _, _, _, _,
  110, -99999, -99999, 235, 230, 200, 220, 235, 235, 240, 235, 235, _, _, _, 
    _, _, _, _, _, _, _,
  260, -99999, 180, 265, 245, 235, 230, 225, 230, 235, 240, 230, _, _, _, _, 
    _, _, _, _, _, _,
  300, -99999, -99999, -99999, 140, 210, 220, 215, 220, 235, 225, 255, _, _, 
    _, _, _, _, _, _, _, _,
  140, -99999, -99999, 155, 200, 210, 210, 215, 215, 215, 220, 235, _, _, _, 
    _, _, _, _, _, _, _,
  0, -99999, 180, 330, 60, 50, 40, 40, 25, 340, 310, 250, _, _, _, _, _, _, 
    _, _, _, _,
  200, -99999, 225, 245, 250, 280, 290, 265, 270, 265, 290, 280, _, _, _, _, 
    _, _, _, _, _, _,
  290, -99999, 310, 275, 265, 270, 265, 255, 255, 255, 260, 255, _, _, _, _, 
    _, _, _, _, _, _,
  340, -99999, -99999, 20, 285, 245, 240, 250, 240, 240, 245, 265, _, _, _, 
    _, _, _, _, _, _, _,
  210, -99999, -99999, 160, 115, 225, 220, 230, 230, 235, 240, 245, _, _, _, 
    _, _, _, _, _, _, _,
  0, 350, 345, 30, 360, 25, 20, 20, 25, 15, 5, 340, _, _, _, _, _, _, _, _, 
    _, _,
  220, -99999, 260, 275, 295, 270, 260, 270, 275, 280, 260, 285, _, _, _, _, 
    _, _, _, _, _, _,
  0, 0, 140, 130, 90, 95, 335, 280, 190, 245, 275, 310, _, _, _, _, _, _, _, 
    _, _, _,
  160, 110, 290, 200, 120, 145, 50, 20, 355, 5, 20, 45, _, _, _, _, _, _, _, 
    _, _, _,
  60, 60, 75, 90, 125, 165, 60, 285, 240, 250, 280, 305, _, _, _, _, _, _, _, 
    _, _, _,
  40, 25, 45, 60, 45, 20, 20, 5, 25, 25, 5, 30, _, _, _, _, _, _, _, _, _, _,
  90, 135, 190, 260, 315, 310, 300, 310, 320, 315, 305, 280, _, _, _, _, _, 
    _, _, _, _, _,
  230, 265, 280, 285, 310, 320, 325, 325, 320, 305, 290, 255, _, _, _, _, _, 
    _, _, _, _, _,
  340, -99999, 345, 330, 290, 280, 275, 270, 265, 265, 265, 270, _, _, _, _, 
    _, _, _, _, _, _,
  330, -99999, 350, 335, 310, 295, 290, 285, 275, 280, 285, 270, _, _, _, _, 
    _, _, _, _, _, _,
  120, 135, 145, 135, 165, 270, 260, 270, 250, 240, 190, 185, _, _, _, _, _, 
    _, _, _, _, _,
  280, 320, 55, 70, 70, 75, 70, 75, 75, 75, 70, 55, _, _, _, _, _, _, _, _, 
    _, _,
  60, 110, 350, 340, 325, 335, 320, 320, 315, 320, 315, 320, _, _, _, _, _, 
    _, _, _, _, _,
  0, 320, 330, 330, 320, 315, 315, 310, 310, 310, 315, 320, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  290, 310, 310, 310, 320, 320, 315, 315, 325, 315, 325, 340, _, _, _, _, _, 
    _, _, _, _, _,
  0, 200, 245, 230, 235, 245, 255, 255, 250, 260, 275, 275, _, _, _, _, _, _, 
    _, _, _, _,
  110, 95, 360, -99999, -99999, -99999, -99999, 220, 275, 280, 265, 205, _, 
    _, _, _, _, _, _, _, _, _,
  90, -99999, 190, 180, 345, 335, 310, 325, 315, 330, 315, 295, _, _, _, _, 
    _, _, _, _, _, _,
  350, 10, 10, 355, 320, 280, 275, 250, 250, 255, 265, 265, _, _, _, _, _, _, 
    _, _, _, _,
  230, 285, 35, 50, 50, 60, 45, 45, 55, 40, 60, 55, _, _, _, _, _, _, _, _, 
    _, _,
  310, 340, 335, 335, 325, 355, 360, 360, 10, 20, 30, 85, _, _, _, _, _, _, 
    _, _, _, _,
  110, 115, 185, 100, 75, 140, 160, 155, 130, 85, 70, 30, _, _, _, _, _, _, 
    _, _, _, _,
  245, 250, 330, 330, 335, 350, 350, 350, 355, 355, 355, 355, _, _, _, _, _, 
    _, _, _, _, _,
  30, -99999, 45, 65, 325, 295, 285, 275, 275, 285, 280, 270, _, _, _, _, _, 
    _, _, _, _, _,
  0, 80, 75, 80, 120, 100, 270, 270, 310, 265, 290, 295, _, _, _, _, _, _, _, 
    _, _, _,
  260, -99999, 290, 230, 215, 215, 225, 220, 230, 235, -99999, -99999, _, _, 
    _, _, _, _, _, _, _, _,
  10, 30, -99999, 100, 155, -99999, -99999, -99999, -99999, -99999, 275, 285, 
    _, _, _, _, _, _, _, _, _, _,
  10, 50, 125, 100, 65, 115, 85, 110, 145, 145, -99999, -99999, _, _, _, _, 
    _, _, _, _, _, _,
  310, -99999, -99999, -99999, -99999, -99999, 250, 250, 235, 235, -99999, 
    -99999, _, _, _, _, _, _, _, _, _, _,
  210, -99999, -99999, 280, 280, 230, 225, 225, 225, 225, 235, 215, _, _, _, 
    _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 0, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 0, _, _, _, _, _, _, _, _, _,
  30, 35, 70, 115, 175, 120, 250, 240, 195, 325, 310, 240, _, _, _, _, _, _, 
    _, _, _, _ ;

 wsMan =
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 1.466015e+13, _, _, _, _, _, _, _, _, _,
  3, 3.6, -99999, 8.2, 8.7, 2.5, 3, 0.5, 14.9, 30.8, 25.7, 12.8, _, _, _, _, 
    _, _, _, _, _, _,
  3, 5.1, 6.1, 5.6, 6.1, 8.2, 11.3, 12.8, 9.7, 6.1, 6.1, 3, _, _, _, _, _, _, 
    _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 1.466015e+13, _, _, _, _, _, _, _, _, _,
  4.1, -99999, 3.6, 2, 9.7, 9.7, 16.4, 22.6, 28.3, 27.2, 23.1, 21.6, 
    1.466015e+13, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 1.466015e+13, _, _, _, _, _, _, _, _, _,
  2, 1.5, 1, 2.5, 1.5, 9.2, 6.6, 6.1, 9.2, 6.1, 15.4, 12.8, _, _, _, _, _, _, 
    _, _, _, _,
  3.6, -99999, 4.1, 2, 7.2, 11.8, 16.9, 21.6, 22.6, 22.6, 16.4, 9.7, _, _, _, 
    _, _, _, _, _, _, _,
  3, 4.6, 7.2, 8.7, 12.8, 22.6, 37, 53, 46.3, 30.8, 17.5, 9.7, _, _, _, _, _, 
    _, _, _, _, _,
  6.6, -99999, -99999, 11.3, 12.3, 18.5, 21.1, 24.7, 28.3, 39.1, 14.9, 9.2, 
    _, _, _, _, _, _, _, _, _, _,
  10.2, 12.3, 15.4, 6.1, 9.2, 12.3, 15.4, 17.5, 21.6, 28.8, 13.8, 6.6, _, _, 
    _, _, _, _, _, _, _, _,
  2, 1.5, 2.5, 4.1, 6.6, 14.9, 14.9, 19, 23.1, 24.7, 15.9, 6.1, _, _, _, _, 
    _, _, _, _, _, _,
  5.6, 2, 3, 5.1, 7.2, 13.3, 14.9, 16.4, 17.5, 21.1, 14.4, 5.6, _, _, _, _, 
    _, _, _, _, _, _,
  4.1, 4.1, 6.1, 9.2, 12.3, 11.3, 12.8, 13.3, 10.8, 15.4, 14.4, 5.1, _, _, _, 
    _, _, _, _, _, _, _,
  1, 1, 2.5, 1.5, 3, 1.5, 1.5, 1, 6.6, 14.9, 28.3, 5.6, _, _, _, _, _, _, _, 
    _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 1.466015e+13, _, _, _, _, _, _, _, _, _,
  2.5, 7.7, 9.2, 10.2, 12.3, 16.9, 28.3, 33.4, 27.7, 22.1, 14.4, 7.7, _, _, 
    _, _, _, _, _, _, _, _,
  3, 5.6, 2.5, 4.6, 8.7, 20.5, 26.2, 35, 36, 41.1, 21.1, 9.2, _, _, _, _, _, 
    _, _, _, _, _,
  1, 1.5, 1, 3.6, 7.7, 23.1, 35.5, 42.2, 45.3, 42.7, 22.1, 7.7, _, _, _, _, 
    _, _, _, _, _, _,
  0.5, 0.5, 2, 3, 11.3, 19.5, 24.1, 31.4, 30.8, 21.1, 12.3, 9.7, _, _, _, _, 
    _, _, _, _, _, _,
  1, 3, 3, 5.6, 9.7, 23.6, 26.2, 31.9, 43.2, 35.5, 20.5, 10.8, _, _, _, _, _, 
    _, _, _, _, _,
  1, 2.5, 2, 2, 10.8, 23.1, 28.8, 33.9, 38, 38.6, 21.1, 8.7, _, _, _, _, _, 
    _, _, _, _, _,
  2.5, 4.6, 4.1, 3.6, 9.2, 23.6, 25.7, 34.4, 32.9, 38, 20, 10.8, _, _, _, _, 
    _, _, _, _, _, _,
  1.5, -99999, 1.5, 4.1, 6.1, 6.6, 6.6, 9.7, 8.7, 10.2, 8.7, 5.1, _, _, _, _, 
    _, _, _, _, _, _,
  3.6, 4.1, 4.6, 2.5, 3, 10.8, 7.2, 10.2, 9.2, 10.8, 15.9, 12.8, _, _, _, _, 
    _, _, _, _, _, _,
  2, 3.6, 2.5, 5.6, 6.1, 3, 3.6, 7.7, 9.7, 6.1, 6.6, 7.2, _, _, _, _, _, _, 
    _, _, _, _,
  4.6, -99999, -99999, -99999, 2, 19.5, 29.3, 35.5, 42.2, 42.2, 25.7, 9.2, _, 
    _, _, _, _, _, _, _, _, _,
  2, -99999, 9.2, 9.7, 10.2, 19.5, 35, 36, 42.7, 48.3, 31.4, 12.8, _, _, _, 
    _, _, _, _, _, _, _,
  1.5, 3, 6.6, 6.6, 7.2, 6.1, 2, 9.2, 14.4, 20.5, 19.5, 18.5, _, _, _, _, _, 
    _, _, _, _, _,
  4.6, 6.1, 13.8, 13.3, 14.4, 28.3, 33.4, 47.3, 44.2, 32.9, 21.1, 10.8, _, _, 
    _, _, _, _, _, _, _, _,
  12.3, 12.3, 11.3, 11.8, 12.8, 9.7, 9.2, 9.7, 8.2, 6.1, 6.1, 6.1, _, _, _, 
    _, _, _, _, _, _, _,
  1, 5.1, 7.7, 8.2, 7.7, 3, 3.6, 6.1, 3.6, 7.7, 11.3, 8.7, _, _, _, _, _, _, 
    _, _, _, _,
  0, 4.1, 7.7, 7.2, 5.6, 2.5, 6.6, 7.7, 7.2, 8.7, 10.8, 5.1, _, _, _, _, _, 
    _, _, _, _, _,
  2, 7.7, 8.7, 4.1, 6.1, 4.6, 4.1, 7.7, 13.3, 15.4, 12.8, 8.2, _, _, _, _, _, 
    _, _, _, _, _,
  0, -99999, 5.6, 5.1, 7.2, 4.6, 7.2, 7.2, 12.8, 17.5, 20, 6.1, _, _, _, _, 
    _, _, _, _, _, _,
  2, 2, 11.8, 11.8, 7.2, 7.2, 9.2, 9.2, 5.6, 5.1, 4.6, 7.2, _, _, _, _, _, _, 
    _, _, _, _,
  7.2, 6.6, 5.1, 5.1, 5.6, 6.1, 10.8, 16.9, 20.5, 30.3, 12.3, 12.3, _, _, _, 
    _, _, _, _, _, _, _,
  4.6, -99999, 14.9, 13.3, 11.8, 11.8, 9.7, 12.8, 13.8, 16.4, 22.1, 7.7, _, 
    _, _, _, _, _, _, _, _, _,
  1.5, 2.5, 6.6, 4.6, 5.1, 13.8, 15.4, 19.5, 25.7, 34.4, 17.5, 12.8, _, _, _, 
    _, _, _, _, _, _, _,
  1, -99999, 8.7, 8.7, 13.8, 9.7, 14.9, 13.8, 22.1, 27.2, 20, 6.6, _, _, _, 
    _, _, _, _, _, _, _,
  4.1, -99999, 16.4, 20, 14.9, 19, 21.1, 17.5, 20.5, 28.3, 20, 10.8, _, _, _, 
    _, _, _, _, _, _, _,
  0, -99999, 3, 3.6, 9.2, 15.4, 23.6, 30.3, 35, 35, 22.6, 13.3, _, _, _, _, 
    _, _, _, _, _, _,
  1.5, 2.5, 4.1, 1.5, 3.6, 14.4, 19, 20.5, 23.1, 28.8, 19.5, 18.5, _, _, _, 
    _, _, _, _, _, _, _,
  2.5, 4.1, 8.7, 8.7, 5.1, 20, 18, 22.1, 21.1, 27.7, 20.5, 14.4, _, _, _, _, 
    _, _, _, _, _, _,
  3.6, -99999, 18.5, 11.8, 14.4, 15.4, 13.3, 16.9, 13.8, 19.5, 15.4, 10.8, _, 
    _, _, _, _, _, _, _, _, _,
  0.5, 3, 4.6, 4.1, 1.5, 4.6, 4.1, 9.7, 14.9, 10.8, 7.2, 8.2, _, _, _, _, _, 
    _, _, _, _, _,
  4.1, -99999, 13.3, 9.7, 12.8, 3, 4.1, 4.6, 5.1, 6.1, 15.4, 13.8, _, _, _, 
    _, _, _, _, _, _, _,
  4.6, -99999, -99999, 13.8, 1.5, 1.5, 8.2, 12.8, 16.9, 20, 20.5, 13.3, _, _, 
    _, _, _, _, _, _, _, _,
  4.6, -99999, -99999, 13.8, 3.6, 6.1, 10.2, 11.8, 12.8, 17.5, 22.1, 14.4, _, 
    _, _, _, _, _, _, _, _, _,
  2.5, -99999, 15.9, 12.3, 2.5, 5.1, 4.6, 5.1, -99999, -99999, 6.1, 4.6, _, 
    _, _, _, _, _, _, _, _, _,
  5.1, -99999, 20.5, 11.3, 9.7, 4.6, 8.2, 8.2, 8.7, 10.8, 14.9, 10.2, _, _, 
    _, _, _, _, _, _, _, _,
  5.6, -99999, -99999, 15.9, 13.3, 9.7, 10.8, 16.4, 13.8, 14.9, 20.5, 16.9, 
    _, _, _, _, _, _, _, _, _, _,
  3.6, -99999, -99999, 6.6, 1.5, 12.3, 17.5, 18.5, 17.5, 24.1, 26.7, 15.9, _, 
    _, _, _, _, _, _, _, _, _,
  2.5, -99999, -99999, -99999, 4.1, 19.5, 17.5, 17.5, 23.6, 25.7, 27.7, 21.6, 
    _, _, _, _, _, _, _, _, _, _,
  2.5, -99999, -99999, -99999, 14.4, 21.6, 17.5, 21.6, 27.7, 33.4, 33.9, 
    14.4, _, _, _, _, _, _, _, _, _, _,
  1.5, -99999, -99999, 3.6, 13.3, 19, 30.3, 38.6, 43.2, 40.1, 21.6, 11.3, _, 
    _, _, _, _, _, _, _, _, _,
  2.5, -99999, 20, 20, 7.7, 5.6, 4.1, 6.1, 8.7, 6.6, 8.7, 5.6, _, _, _, _, _, 
    _, _, _, _, _,
  4.6, -99999, -99999, 22.1, 18, 10.8, 14.9, 18.5, 20, 21.1, 22.6, 9.7, _, _, 
    _, _, _, _, _, _, _, _,
  3, -99999, -99999, -99999, 3, 21.1, 17.5, 19.5, 25.7, 34.4, 25.2, 15.4, _, 
    _, _, _, _, _, _, _, _, _,
  5.1, -99999, -99999, -99999, 7.7, 19.5, 24.7, 28.3, 30.3, 33.4, 27.2, 19, 
    _, _, _, _, _, _, _, _, _, _,
  3.6, 4.1, 4.1, 2.5, 5.1, 5.6, 5.1, 18, 15.9, 14.9, 9.7, 12.8, _, _, _, _, 
    _, _, _, _, _, _,
  2.5, -99999, -99999, 4.1, 12.3, 19.5, 21.1, 28.3, 30.8, 27.2, 22.6, 9.2, _, 
    _, _, _, _, _, _, _, _, _,
  3.6, -99999, -99999, 15.4, 6.1, 23.6, 25.7, 24.7, 26.7, 28.3, 21.6, 14.9, 
    _, _, _, _, _, _, _, _, _, _,
  1, -99999, -99999, -99999, 2.5, 12.8, 22.1, 33.4, 33.9, 29.8, 22.1, 11.8, 
    _, _, _, _, _, _, _, _, _, _,
  3, -99999, 12.8, 15.9, 14.9, 33.4, 32.9, 32.4, 30.3, 28.3, 34.4, 12.8, _, 
    _, _, _, _, _, _, _, _, _,
  8.7, -99999, 18.5, 11.8, 12.3, 27.7, 36, 39.6, 46.3, 48.9, 30.3, 15.4, _, 
    _, _, _, _, _, _, _, _, _,
  2, -99999, -99999, 2.5, 4.6, 11.3, 16.4, 21.6, 24.7, 14.9, 15.9, 10.8, _, 
    _, _, _, _, _, _, _, _, _,
  4.6, -99999, 13.8, 12.3, 14.4, 26.2, 29.3, 44.7, 46.8, 45.3, 32.4, 14.4, _, 
    _, _, _, _, _, _, _, _, _,
  1.5, -99999, 2.5, 2.5, 1.5, 8.2, 12.8, 36, 43.7, 40.6, 23.1, 12.8, _, _, _, 
    _, _, _, _, _, _, _,
  2, -99999, 2.5, 2, 1.5, 3.6, 1.5, 6.1, 7.2, 5.1, 6.1, 6.6, _, _, _, _, _, 
    _, _, _, _, _,
  4.6, 5.1, 6.6, 3.6, 1.5, 5.6, 5.6, 6.6, 7.2, 4.6, 15.9, 9.2, _, _, _, _, _, 
    _, _, _, _, _,
  2.5, 8.7, 8.2, 6.6, 6.6, 12.3, 15.9, 14.4, 10.8, 8.7, 7.7, 6.1, _, _, _, _, 
    _, _, _, _, _, _,
  0, 3.6, 3, 5.6, 8.7, 12.8, 23.1, 26.2, 29.8, 23.1, 19, 11.8, _, _, _, _, _, 
    _, _, _, _, _,
  2.5, -99999, 12.3, 12.8, 12.8, 19.5, 22.1, 29.8, 44.2, 50.9, 26.2, 16.4, _, 
    _, _, _, _, _, _, _, _, _,
  2, 1.5, 8.7, 12.3, 14.4, 26.2, 28.3, 32.4, 25.2, 25.7, 20, 11.8, _, _, _, 
    _, _, _, _, _, _, _,
  5.1, 5.1, 12.8, 13.8, 15.4, 22.6, 28.3, 29.3, 36.5, 21.6, 14.4, 4.6, _, _, 
    _, _, _, _, _, _, _, _,
  7.7, -99999, 6.6, 12.3, 21.6, 32.4, 36, 37.5, 31.4, 23.6, 15.9, 5.1, _, _, 
    _, _, _, _, _, _, _, _,
  2.5, 3.6, 3, 1.5, 8.2, 8.2, 13.3, 18, 23.1, 29.3, 22.1, 8.7, _, _, _, _, _, 
    _, _, _, _, _,
  3.6, 6.6, 10.2, 9.2, 4.6, 2.5, 5.1, 3.6, 10.8, 20.5, 20.5, 9.7, _, _, _, _, 
    _, _, _, _, _, _,
  1.5, 4.6, 1, 3.6, 4.6, 0.5, 4.6, 4.6, 7.2, 7.2, 7.7, 4.6, _, _, _, _, _, _, 
    _, _, _, _,
  2.5, 6.1, 3.6, 1, 1, 4.6, 3.6, 6.6, 9.7, 14.9, 11.3, 7.2, _, _, _, _, _, _, 
    _, _, _, _,
  0, 1.5, 1, -99999, -99999, 3.6, 2, 5.1, 7.7, 7.7, 8.2, 4.6, _, _, _, _, _, 
    _, _, _, _, _,
  1, -99999, 4.6, 3, 2.5, 2.5, 5.6, 5.6, 9.7, 11.3, 8.2, 6.6, _, _, _, _, _, 
    _, _, _, _, _,
  1, 5.1, 7.7, 9.2, 7.7, 5.6, -99999, -99999, -99999, -99999, -99999, -99999, 
    _, _, _, _, _, _, _, _, _, _,
  2, 5.1, 10.8, 7.7, 11.3, 4.1, 7.7, 3, 0.5, 4.6, 4.1, -99999, _, _, _, _, _, 
    _, _, _, _, _,
  0, -99999, 5.1, 8.2, 9.2, 5.1, 7.7, 9.2, 13.3, 16.4, 20, 7.2, _, _, _, _, 
    _, _, _, _, _, _,
  0.5, 3.6, 8.7, 4.6, 6.1, 11.8, 16.4, 19.5, 22.6, 25.7, 17.5, 15.4, _, _, _, 
    _, _, _, _, _, _, _,
  3, -99999, -99999, 10.8, 12.8, 12.8, 16.9, 27.7, 29.8, 38.6, 21.1, 11.3, _, 
    _, _, _, _, _, _, _, _, _,
  3, 6.6, 10.2, 9.2, 4.6, 11.8, 16.4, 26.2, 29.8, 30.8, 31.4, 15.9, _, _, _, 
    _, _, _, _, _, _, _,
  4.6, 7.7, 10.8, 9.7, 3.6, 4.6, 7.7, 10.2, 14.9, 24.7, 27.2, 18, _, _, _, _, 
    _, _, _, _, _, _,
  2.5, 6.6, 11.8, 10.8, 3.6, 5.1, 7.2, 7.2, 12.3, 10.8, 25.2, 15.9, _, _, _, 
    _, _, _, _, _, _, _,
  2.5, -99999, -99999, 3.6, 13.3, 23.1, 18.5, 21.6, 29.3, 35.5, 25.7, 15.4, 
    _, _, _, _, _, _, _, _, _, _,
  2, -99999, 1.5, 6.1, 15.4, 22.6, 32.4, 35.5, 40.6, 43.7, 36, 13.3, _, _, _, 
    _, _, _, _, _, _, _,
  1.5, -99999, -99999, -99999, 3.6, 10.2, 11.3, 18, 18, 19, 11.8, 8.2, _, _, 
    _, _, _, _, _, _, _, _,
  2, -99999, -99999, 4.6, 9.2, 19, 27.2, 37, 40.1, 38, 23.6, 15.4, _, _, _, 
    _, _, _, _, _, _, _,
  0, -99999, 2, 1, 2, 8.7, 13.3, 14.9, 10.2, 4.6, 4.1, 7.2, _, _, _, _, _, _, 
    _, _, _, _,
  5.1, -99999, 26.2, 22.1, 20, 30.8, 30.8, 25.2, 27.2, 41.1, 37, 13.8, _, _, 
    _, _, _, _, _, _, _, _,
  2, -99999, 9.7, 12.3, 27.7, 37.5, 37, 40.1, 47.3, 53.5, 46.3, 18.5, _, _, 
    _, _, _, _, _, _, _, _,
  2.5, -99999, -99999, 8.2, 4.6, 22.6, 27.2, 34.4, 35.5, 39.6, 30.8, 14.9, _, 
    _, _, _, _, _, _, _, _, _,
  3.6, -99999, -99999, 5.1, 7.2, 9.7, 8.2, 22.6, 31.9, 23.6, 19, 12.8, _, _, 
    _, _, _, _, _, _, _, _,
  0, 1, 4.1, 7.2, 5.6, 7.2, 16.9, 24.1, 30.3, 23.6, 11.8, 7.2, _, _, _, _, _, 
    _, _, _, _, _,
  6.1, -99999, 16.4, 10.8, 13.3, 20.5, 26.2, 23.1, 22.6, 25.2, 21.1, 14.9, _, 
    _, _, _, _, _, _, _, _, _,
  0, 0, 2, 1.5, 3, 2.5, 5.1, 5.6, 6.6, 12.3, 16.4, 14.9, _, _, _, _, _, _, _, 
    _, _, _,
  2, 1.5, 1, 3, 4.1, 3, 2, 12.8, 16.9, 15.4, 33.4, 18, _, _, _, _, _, _, _, 
    _, _, _,
  4.6, 4.6, 3.6, 3, 4.1, 2.5, 3, 6.1, 11.8, 12.3, 15.9, 19.5, _, _, _, _, _, 
    _, _, _, _, _,
  1, 1.5, 2.5, 4.6, 5.1, 10.8, 12.3, 8.2, 9.2, 8.7, 7.7, 5.6, _, _, _, _, _, 
    _, _, _, _, _,
  1, 2.5, 7.2, 6.6, 13.3, 19, 25.2, 34.4, 42.7, 36.5, 23.1, 11.3, _, _, _, _, 
    _, _, _, _, _, _,
  4.1, 6.1, 8.7, 12.3, 15.9, 29.8, 35, 40.1, 36.5, 23.6, 10.2, 6.1, _, _, _, 
    _, _, _, _, _, _, _,
  7.7, -99999, 10.2, 11.8, 17.5, 26.7, 30.3, 37, 38.6, 36, 31.9, 18, _, _, _, 
    _, _, _, _, _, _, _,
  5.1, -99999, 7.2, 14.9, 21.1, 29.8, 35.5, 40.1, 36, 31.9, 24.1, 13.8, _, _, 
    _, _, _, _, _, _, _, _,
  3.6, 6.1, 7.7, 10.2, 7.2, 10.8, 15.9, 18, 10.2, 8.2, 7.2, 3.6, _, _, _, _, 
    _, _, _, _, _, _,
  3, 2.5, 3.6, 7.7, 8.7, 9.7, 12.8, 13.3, 10.2, 8.2, 6.1, 5.1, _, _, _, _, _, 
    _, _, _, _, _,
  1, 2.5, 3, 8.2, 12.3, 24.7, 22.6, 17.5, 17.5, 14.9, 14.9, 8.7, _, _, _, _, 
    _, _, _, _, _, _,
  0, 7.7, 11.3, 12.8, 12.3, 10.2, 15.9, 15.4, 14.4, 14.9, 9.2, 7.2, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.6, 12.8, 20, 21.1, 13.8, 15.4, 26.7, 26.7, 21.1, 14.4, 11.3, 9.7, _, _, 
    _, _, _, _, _, _, _, _,
  0, 1, 11.3, 18, 27.2, 25.7, 25.7, 34.4, 42.2, 45.3, 27.2, 13.3, _, _, _, _, 
    _, _, _, _, _, _,
  2.5, 2, 5.6, -99999, -99999, -99999, -99999, 4.1, 10.2, 18, 20.5, 3.6, _, 
    _, _, _, _, _, _, _, _, _,
  0.5, -99999, 5.6, 2.5, 4.6, 3.6, 6.1, 10.8, 8.2, 8.2, 7.2, 6.6, _, _, _, _, 
    _, _, _, _, _, _,
  3.6, 7.7, 10.2, 16.9, 12.8, 18, 21.1, 39.1, 50.4, 30.8, 18.5, 8.2, _, _, _, 
    _, _, _, _, _, _, _,
  1, 3.6, 6.6, 9.2, 8.7, 10.8, 8.7, 13.8, 9.7, 4.6, 3.6, 2, _, _, _, _, _, _, 
    _, _, _, _,
  3, 6.1, 7.2, 7.7, 4.6, 4.6, 8.7, 11.8, 9.7, 9.2, 7.2, 3.6, _, _, _, _, _, 
    _, _, _, _, _,
  4.1, 5.1, 2, 2, 6.1, 5.1, 11.8, 14.9, 8.2, 15.9, 14.9, 8.7, _, _, _, _, _, 
    _, _, _, _, _,
  2.5, 2, 4.1, 5.6, 6.1, 21.6, 22.6, 28.8, 30.8, 39.1, 12.3, 8.7, _, _, _, _, 
    _, _, _, _, _, _,
  1.5, -99999, 4.1, 9.7, 9.2, 11.8, 11.3, 18.5, 24.7, 15.4, 12.8, 10.2, _, _, 
    _, _, _, _, _, _, _, _,
  0, 6.6, 9.2, 9.7, 7.2, 3, 7.2, 14.9, 21.6, 19.5, 23.1, 11.8, _, _, _, _, _, 
    _, _, _, _, _,
  0.5, -99999, 8.7, 8.2, 11.3, 22.6, 25.7, 31.9, 37, 42.7, -99999, -99999, _, 
    _, _, _, _, _, _, _, _, _,
  4.1, 3.6, -99999, 9.2, 2.5, -99999, -99999, -99999, -99999, -99999, 26.2, 
    15.4, _, _, _, _, _, _, _, _, _, _,
  1.5, 2.5, 4.6, 5.1, 5.1, 3.6, 4.1, 3.6, 2.5, 4.1, -99999, -99999, _, _, _, 
    _, _, _, _, _, _, _,
  5.1, -99999, -99999, -99999, -99999, -99999, 25.2, 36.5, 41.1, 39.6, 
    -99999, -99999, _, _, _, _, _, _, _, _, _, _,
  7.2, -99999, -99999, 10.2, 6.6, 18, 24.1, 31.4, 42.2, 37, 26.7, 12.8, _, _, 
    _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 1.466015e+13, _, _, _, _, _, _, _, _, _,
  -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, -99999, 
    -99999, -99999, -99999, 1.466015e+13, _, _, _, _, _, _, _, _, _,
  1.5, 1.5, 4.1, 7.2, 1, 7.2, 13.8, 11.8, 5.1, 7.2, 5.1, 2.5, _, _, _, _, _, 
    _, _, _, _, _ ;

 prSigT =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1021, 904, 889, 835, 780, 770, 759, 695, 676, 589, 481, 255, 157, 100, 
    10000, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1029, 1018, 768, 625, 574, 500, 324, 211, 150, 100, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1005, 1004, 939, 937, 922, 917, 916, 915, 897, 875, 873, 867, 850, 819, 
    791, 770, 769, 767, 766, 763, 762, 739, 707, 676, 524, 385, 365, 351, 
    308, 290, 238, 233, 212, 210, 204, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  979, 942, 874, 762, 636, 614, 610, 594, 586, 536, 520, 508, 457, 453, 416, 
    393, 363, 330, 306, 278, 262, 218, 189, 173, 146, 119, 111, 101, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1002, 971, 910, 799, 792, 782, 732, 690, 653, 629, 610, 595, 564, 537, 422, 
    384, 337, 261, 239, 212, 200, 131, 100, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1021, 957, 887, 812, 740, 580, 500, 231, 188, 164, 159, 124, 100, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  944, 938, 914, 911, 885, 883, 866, 850, 792, 643, 400, 178, 162, 111, 102, 
    100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  997, 981, 864, 861, 840, 775, 702, 700, 687, 611, 572, 545, 500, 436, 374, 
    345, 293, 178, 155, 139, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1000, 956, 925, 871, 835, 826, 776, 617, 611, 604, 589, 583, 560, 555, 535, 
    475, 318, 292, 175, 150, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  977, 898, 887, 878, 776, 768, 754, 714, 686, 680, 570, 552, 548, 538, 496, 
    453, 434, 423, 391, 378, 324, 300, 295, 270, 187, 103, 100, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  984, 887, 776, 751, 737, 727, 714, 669, 598, 574, 565, 459, 450, 440, 434, 
    428, 400, 364, 354, 337, 300, 141, 100, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1032, 1015, 850, 808, 736, 730, 724, 695, 682, 630, 594, 482, 472, 449, 
    432, 330, 277, 193, 171, 156, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1017, 850, 837, 826, 811, 802, 711, 682, 667, 657, 649, 640, 611, 588, 526, 
    458, 421, 337, 321, 180, 168, 137, 108, 100, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1006, 988, 900, 850, 815, 760, 757, 750, 718, 700, 675, 661, 654, 645, 641, 
    617, 440, 427, 380, 330, 208, 171, 119, 100, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  987, 925, 770, 700, 653, 646, 621, 606, 595, 588, 577, 557, 543, 527, 517, 
    509, 485, 470, 446, 394, 375, 326, 280, 221, 184, 152, 100, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1025, 1009, 995, 896, 862, 840, 785, 765, 756, 741, 712, 619, 606, 500, 
    450, 400, 318, 259, 188, 170, 150, 111, 100, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  951, 946, 895, 864, 747, 709, 687, 671, 500, 466, 282, 195, 165, 118, 100, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1008, 997, 958, 925, 850, 700, 518, 458, 375, 338, 266, 183, 157, 100, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  996, 925, 860, 831, 774, 684, 645, 580, 575, 539, 523, 496, 490, 488, 484, 
    483, 480, 473, 469, 462, 438, 400, 393, 381, 374, 370, 355, 349, 338, 
    325, 303, 293, 279, 269, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  890, 734, 678, 576, 414, 375, 339, 312, 264, 245, 150, 108, 100, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1021, 1005, 925, 907, 900, 880, 811, 799, 772, 767, 729, 724, 721, 714, 
    700, 657, 595, 581, 553, 382, 211, 173, 154, 145, 131, 100, 10000, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  799, 712, 681, 669, 621, 602, 488, 476, 450, 431, 400, 382, 342, 222, 191, 
    185, 123, 112, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  955, 908, 837, 819, 753, 700, 667, 650, 642, 635, 623, 618, 616, 604, 595, 
    579, 573, 564, 562, 560, 528, 524, 519, 500, 495, 422, 414, 400, 260, 
    188, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1007, 798, 790, 781, 729, 710, 663, 659, 651, 633, 606, 572, 550, 500, 489, 
    451, 445, 434, 429, 413, 404, 396, 387, 360, 354, 349, 330, 316, 300, 
    287, 270, 184, 129, 106, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1004, 951, 933, 881, 808, 774, 721, 678, 594, 372, 290, 259, 220, 197, 182, 
    174, 140, 133, 110, 101, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  994, 982, 934, 848, 836, 818, 812, 787, 769, 763, 751, 709, 627, 559, 533, 
    505, 413, 341, 301, 279, 258, 251, 236, 221, 213, 188, 173, 162, 148, 
    139, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1021, 1017, 951, 906, 850, 798, 776, 773, 760, 756, 753, 700, 641, 636, 
    623, 575, 500, 206, 105, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1000, 981, 947, 902, 891, 883, 873, 863, 839, 821, 744, 725, 717, 695, 655, 
    631, 553, 533, 530, 520, 516, 479, 472, 437, 425, 404, 395, 368, 177, 
    141, 125, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1014, 984, 975, 969, 962, 943, 804, 663, 631, 623, 589, 574, 540, 528, 520, 
    506, 477, 462, 443, 367, 339, 326, 300, 169, 133, 100, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  955, 805, 632, 628, 623, 611, 577, 568, 517, 511, 493, 474, 422, 400, 279, 
    263, 239, 176, 142, 138, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  985, 960, 886, 822, 714, 695, 688, 683, 679, 648, 636, 611, 600, 506, 496, 
    460, 437, 417, 393, 372, 361, 330, 250, 150, 126, 119, 100, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1012, 826, 770, 708, 671, 665, 655, 630, 479, 449, 331, 316, 176, 164, 151, 
    134, 132, 129, 123, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  960, 944, 716, 711, 704, 626, 591, 538, 532, 520, 448, 345, 226, 178, 139, 
    100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  996, 991, 980, 942, 865, 794, 659, 629, 539, 474, 400, 388, 313, 257, 193, 
    174, 173, 155, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  962, 951, 916, 824, 700, 695, 658, 643, 613, 598, 526, 521, 500, 480, 450, 
    323, 200, 142, 106, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  944, 933, 910, 834, 757, 718, 713, 686, 649, 627, 575, 536, 440, 344, 188, 
    171, 162, 158, 138, 131, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  992, 966, 823, 777, 668, 653, 484, 466, 417, 400, 384, 329, 225, 192, 182, 
    100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1010, 986, 812, 806, 779, 604, 598, 596, 592, 549, 529, 481, 475, 409, 314, 
    260, 225, 181, 168, 117, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1015, 1004, 992, 850, 817, 633, 578, 500, 250, 194, 188, 166, 100, 192, 
    182, 100, 162, 158, 138, 131, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  993, 955, 948, 850, 801, 747, 733, 725, 568, 400, 362, 259, 240, 163, 131, 
    126, 108, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1021, 1012, 967, 902, 894, 876, 864, 829, 740, 670, 657, 638, 632, 573, 
    543, 540, 529, 525, 489, 461, 452, 442, 420, 408, 300, 185, 150, 141, 
    131, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  995, 951, 912, 880, 806, 781, 778, 736, 587, 515, 176, 125, 100, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  879, 867, 802, 758, 752, 742, 731, 723, 700, 598, 537, 339, 167, 100, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  850, 818, 802, 762, 370, 327, 322, 300, 209, 140, 130, 104, 100, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  959, 946, 903, 850, 790, 647, 623, 601, 537, 512, 484, 477, 460, 383, 147, 
    109, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  943, 925, 891, 870, 857, 850, 835, 801, 583, 579, 545, 383, 300, 260, 164, 
    143, 116, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  858, 840, 829, 826, 774, 652, 565, 525, 515, 472, 426, 391, 381, 371, 350, 
    304, 282, 233, 172, 150, 120, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  865, 760, 654, 535, 529, 433, 400, 376, 326, 255, 177, 141, 128, 114, 100, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  826, 755, 726, 695, 599, 486, 474, 471, 464, 435, 400, 343, 300, 289, 274, 
    167, 124, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  771, 651, 642, 613, 586, 546, 475, 469, 464, 375, 319, 311, 300, 274, 190, 
    173, 141, 116, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  800, 729, 604, 438, 421, 407, 400, 216, 164, 100, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  956, 881, 876, 855, 845, 728, 556, 536, 527, 524, 522, 443, 335, 313, 250, 
    200, 139, 127, 117, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  897, 880, 585, 500, 462, 426, 400, 352, 342, 323, 311, 155, 130, 100, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  703, 687, 634, 621, 619, 613, 601, 460, 449, 445, 421, 374, 359, 300, 183, 
    145, 128, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  828, 750, 555, 545, 523, 519, 509, 472, 459, 352, 189, 174, 131, 116, 107, 
    100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  982, 941, 919, 887, 877, 848, 841, 820, 814, 795, 730, 724, 702, 700, 537, 
    349, 270, 250, 215, 176, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  901, 884, 838, 797, 778, 700, 637, 512, 455, 442, 359, 325, 313, 300, 279, 
    250, 183, 143, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  868, 864, 859, 832, 825, 802, 756, 683, 674, 656, 632, 460, 431, 411, 405, 
    400, 357, 278, 243, 231, 200, 155, 114, 100, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  836, 818, 750, 680, 635, 574, 532, 500, 491, 484, 479, 351, 250, 218, 171, 
    100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  913, 897, 820, 734, 662, 647, 633, 607, 581, 556, 542, 533, 526, 508, 500, 
    400, 187, 150, 127, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  885, 872, 799, 753, 729, 700, 670, 651, 639, 600, 576, 532, 483, 435, 409, 
    390, 352, 311, 300, 225, 173, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  907, 900, 896, 888, 868, 681, 596, 559, 500, 460, 430, 316, 247, 200, 175, 
    100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  892, 875, 803, 797, 783, 700, 683, 643, 608, 592, 556, 520, 510, 491, 387, 
    354, 344, 329, 265, 250, 174, 154, 140, 100, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  930, 927, 925, 905, 761, 666, 652, 629, 618, 549, 453, 438, 424, 371, 356, 
    337, 228, 207, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  925, 879, 823, 661, 614, 608, 577, 535, 521, 500, 432, 238, 192, 132, 100, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1000, 890, 836, 829, 799, 783, 748, 739, 715, 684, 651, 636, 626, 621, 616, 
    614, 571, 540, 530, 500, 436, 384, 376, 365, 187, 110, 100, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1011, 1004, 985, 967, 894, 845, 821, 776, 729, 661, 651, 567, 514, 472, 
    426, 405, 321, 306, 275, 238, 227, 223, 203, 142, 100, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1003, 989, 971, 923, 804, 757, 732, 583, 494, 396, 327, 277, 231, 221, 203, 
    189, 173, 157, 133, 114, 107, 104, 100, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  964, 829, 813, 802, 630, 528, 512, 501, 464, 450, 414, 389, 340, 296, 258, 
    213, 188, 182, 171, 147, 144, 135, 110, 100, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1011, 988, 966, 928, 866, 823, 799, 791, 773, 768, 719, 638, 517, 383, 292, 
    248, 213, 198, 166, 141, 135, 115, 100, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  957, 932, 894, 851, 822, 673, 564, 352, 243, 235, 218, 203, 192, 154, 134, 
    125, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  953, 940, 900, 885, 875, 853, 843, 819, 813, 728, 527, 372, 290, 257, 248, 
    239, 229, 201, 183, 158, 155, 146, 133, 110, 100, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1013, 925, 791, 748, 718, 716, 713, 680, 675, 663, 656, 601, 500, 461, 416, 
    386, 333, 315, 215, 157, 146, 142, 130, 115, 100, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1020, 1018, 956, 925, 848, 772, 755, 722, 593, 535, 500, 496, 491, 485, 
    469, 460, 417, 392, 378, 359, 341, 327, 266, 163, 151, 144, 102, 100, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1000, 964, 934, 925, 881, 832, 803, 758, 717, 600, 578, 427, 414, 400, 347, 
    312, 200, 158, 135, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1007, 968, 953, 913, 770, 619, 576, 538, 520, 443, 418, 339, 310, 288, 167, 
    143, 139, 111, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1004, 870, 829, 766, 700, 574, 548, 537, 510, 488, 472, 464, 400, 339, 185, 
    148, 128, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  985, 967, 775, 673, 615, 571, 549, 545, 475, 426, 387, 380, 351, 309, 250, 
    200, 148, 128, 117, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1012, 929, 887, 884, 861, 850, 764, 745, 718, 709, 697, 651, 622, 599, 591, 
    581, 565, 532, 513, 496, 449, 409, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  925, 912, 898, 890, 850, 815, 799, 760, 758, 737, 700, 569, 500, 469, 326, 
    173, 150, 132, 111, 105, 1000, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  939, 932, 907, 850, 662, 628, 605, 598, 590, 532, 434, 313, 300, 250, 204, 
    143, 115, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1006, 992, 982, 968, 960, 939, 869, 850, 824, 682, 574, 451, 391, 383, 353, 
    340, 227, 172, 132, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  950, 857, 844, 828, 797, 743, 682, 629, 601, 515, 482, 474, 419, 369, 209, 
    187, 175, 142, 122, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1000, 925, 884, 786, 744, 736, 733, 717, 658, 630, 602, 588, 572, 552, 544, 
    517, 484, 482, 472, 448, 433, 388, 314, 300, 269, 250, 117, 100, 116, 
    100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1000, 899, 868, 817, 809, 761, 706, 688, 666, 603, 538, 163, 100, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1000, 925, 850, 824, 805, 779, 747, 727, 700, 677, 672, 659, 619, 558, 422, 
    396, 182, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  903, 787, 715, 666, 650, 588, 483, 448, 300, 267, 227, 195, 143, 133, 114, 
    100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  925, 893, 887, 877, 850, 826, 709, 681, 632, 542, 525, 469, 381, 365, 332, 
    316, 200, 175, 135, 105, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  758, 750, 735, 685, 673, 658, 653, 471, 370, 321, 236, 154, 114, 100, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  863, 850, 800, 731, 646, 600, 580, 558, 532, 505, 500, 475, 463, 444, 434, 
    400, 369, 345, 311, 288, 208, 192, 158, 121, 100, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  948, 878, 850, 817, 787, 778, 760, 687, 679, 671, 650, 630, 622, 612, 599, 
    588, 583, 573, 557, 500, 388, 369, 335, 269, 240, 168, 100, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  941, 933, 919, 912, 850, 781, 667, 605, 595, 551, 543, 522, 507, 493, 452, 
    444, 430, 423, 416, 366, 361, 344, 162, 150, 138, 122, 117, 100, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  935, 918, 770, 747, 710, 698, 691, 646, 639, 624, 589, 565, 528, 477, 442, 
    415, 409, 377, 300, 285, 265, 250, 158, 145, 135, 128, 104, 100, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  888, 808, 798, 765, 745, 700, 665, 622, 588, 500, 360, 240, 160, 148, 139, 
    135, 120, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  883, 870, 822, 674, 642, 631, 591, 540, 529, 517, 500, 490, 425, 374, 347, 
    321, 230, 166, 100, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  925, 899, 860, 855, 840, 820, 581, 571, 560, 541, 534, 527, 522, 481, 461, 
    400, 340, 217, 176, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  876, 832, 819, 760, 727, 580, 568, 530, 356, 250, 215, 179, 134, 123, 110, 
    103, 100, 217, 176, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  925, 718, 714, 706, 658, 651, 591, 535, 519, 512, 463, 449, 445, 442, 439, 
    433, 343, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  890, 875, 844, 832, 824, 807, 782, 665, 658, 652, 648, 616, 580, 571, 538, 
    504, 489, 470, 451, 440, 429, 376, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  955, 689, 681, 674, 663, 653, 440, 261, 125, 108, 100, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  1016, 1008, 973, 959, 947, 891, 849, 838, 832, 821, 809, 766, 619, 591, 
    569, 462, 409, 378, 350, 277, 236, 183, 140, 116, 100, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  997, 978, 852, 831, 792, 775, 765, 721, 707, 593, 542, 497, 476, 459, 433, 
    417, 401, 346, 318, 224, 210, 193, 168, 144, 136, 128, 116, 101, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1009, 845, 840, 831, 813, 711, 597, 582, 528, 489, 397, 313, 262, 257, 245, 
    235, 221, 204, 165, 149, 120, 113, 101, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  892, 880, 874, 856, 825, 813, 807, 801, 789, 783, 753, 714, 704, 607, 516, 
    475, 355, 251, 235, 198, 181, 151, 143, 132, 121, 112, 107, 101, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  979, 916, 900, 884, 855, 615, 592, 583, 547, 522, 511, 416, 332, 283, 243, 
    237, 228, 223, 206, 194, 178, 171, 155, 118, 114, 100, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  998, 965, 910, 819, 813, 807, 705, 578, 556, 513, 510, 473, 423, 411, 401, 
    351, 289, 257, 244, 175, 101, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  995, 989, 928, 892, 887, 882, 847, 801, 769, 684, 617, 562, 530, 518, 477, 
    453, 397, 349, 306, 285, 236, 217, 187, 154, 108, 103, 101, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  998, 876, 858, 846, 812, 785, 774, 759, 725, 706, 670, 631, 611, 593, 559, 
    543, 473, 452, 414, 317, 292, 272, 261, 254, 234, 224, 160, 118, 100, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  994, 983, 965, 826, 784, 738, 720, 686, 663, 402, 319, 301, 285, 276, 267, 
    252, 211, 194, 166, 141, 131, 109, 100, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  923, 784, 723, 636, 629, 589, 582, 575, 566, 561, 496, 479, 467, 418, 393, 
    371, 332, 302, 230, 202, 183, 165, 154, 138, 118, 109, 100, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1017, 931, 899, 766, 729, 537, 491, 464, 349, 305, 281, 249, 224, 187, 152, 
    117, 110, 101, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  992, 760, 562, 506, 482, 467, 445, 388, 375, 284, 263, 234, 219, 190, 160, 
    157, 137, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1008, 875, 731, 692, 683, 675, 648, 646, 638, 599, 501, 498, 485, 451, 433, 
    405, 375, 282, 186, 142, 126, 107, 107, 10700, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  961, 953, 915, 789, 562, 539, 518, 508, 497, 475, 427, 375, 346, 326, 304, 
    237, 207, 201, 182, 170, 160, 150, 141, 131, 107, 100, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1020, 993, 915, 848, 820, 749, 719, 505, 347, 287, 275, 251, 231, 219, 191, 
    184, 180, 154, 147, 121, 113, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1008, 976, 951, 938, 884, 847, 748, 721, 653, 560, 441, 304, 273, 247, 230, 
    201, 128, 104, 101, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1015, 870, 864, 840, 815, 810, 782, 694, 631, 594, 554, 467, 389, 257, 155, 
    119, 106, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1017, 951, 945, 935, 898, 872, 862, 711, 699, 682, 632, 597, 590, 574, 531, 
    508, 427, 357, 344, 280, 192, 187, 170, 153, 140, 112, 100, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  917, 876, 761, 756, 753, 709, 649, 628, 581, 546, 528, 498, 485, 364, 247, 
    235, 219, 189, 177, 171, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1016, 982, 847, 789, 777, 760, 729, 711, 700, 640, 630, 614, 599, 549, 540, 
    533, 462, 458, 441, 421, 406, 402, 393, 378, 325, 296, 197, 180, 135, 
    105, 105, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  924, 814, 783, 626, 603, 557, 544, 535, 522, 488, 463, 420, 412, 396, 380, 
    315, 309, 197, 190, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1015, 955, 928, 894, 873, 799, 789, 764, 730, 710, 689, 684, 679, 674, 643, 
    636, 632, 623, 620, 600, 578, 575, 569, 540, 537, 491, 449, 442, 416, 
    410, 394, 384, 384, 38400, 38400, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  1016, 1015, 995, 976, 961, 952, 939, 876, 790, 783, 728, 673, 616, 588, 
    487, 397, 349, 336, 299, 250, 201, 198, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1016, 1012, 941, 918, 905, 897, 834, 798, 786, 779, 649, 529, 483, 402, 
    295, 214, 192, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  930, 923, 895, 820, 757, 571, 542, 401, 288, 181, 155, 100, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1007, 984, 945, 840, 772, 693, 674, 649, 631, 610, 456, 406, 291, 177, 134, 
    118, 106, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 tpSigT =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  296.1, 289.1, 288.9, 284.7, 281.5, 281.1, 282.9, 278.1, 277.5, 273.5, 
    262.2, 226.8, 207.8, 205.4, 205.4, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  272.6, 276.1, 260, 250.4, 247.4, 241.8, 221.6, 229.2, 229.4, 224.2, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  283.9, 283.9, 279.9, 279.9, 280.5, 280.9, 280.7, 280.7, 283.9, 285.7, 
    285.7, 285.1, 283.5, 280.5, 278.5, 276.5, 276.5, 276.3, 276.3, 277.7, 
    277.7, 276.7, 275.3, 273, 257, 241.6, 241.2, 239.2, 228.8, 228.6, 224.2, 
    225.2, 222.6, 222, 222.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  280.9, 278.9, 273.7, 268.8, 258.6, 257.2, 257, 255.8, 255.4, 251.6, 250.4, 
    248.8, 242, 241.4, 237.6, 235, 230, 224.6, 222, 218.6, 217, 222.6, 224.2, 
    223.8, 225.4, 221.6, 223.8, 220.4, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  272.6, 273.1, 270.8, 263.2, 263.4, 263.8, 260.6, 261, 259, 258.6, 257.2, 
    256, 254, 251.6, 237.6, 236, 228.8, 219.2, 224, 222, 224.4, 224.8, 221, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  277.3, 276.9, 273.1, 271, 271.4, 263.4, 256.6, 216.2, 209.8, 213.2, 217, 
    220.2, 219, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  274.5, 275.7, 275.3, 277.1, 281.1, 282.1, 281.3, 280.3, 276.5, 269.4, 
    246.6, 206.2, 212.2, 218.6, 216.8, 216.8, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  279.9, 280.5, 273.7, 275.5, 276.7, 275.9, 272.6, 272.6, 271, 265, 263.8, 
    260.6, 257, 249, 241.2, 236.4, 230.8, 205.8, 213.6, 216, 217.8, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  281.3, 280.3, 280.5, 278.7, 277.9, 277.5, 277.1, 268.2, 268, 267.6, 266.4, 
    266, 263.8, 263.2, 261, 253.8, 232.4, 231.4, 206, 213.8, 216.2, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  295.5, 291.5, 290.9, 290.5, 283.7, 284.1, 283.9, 280.7, 279.3, 278.9, 
    271.6, 270, 269.6, 268.4, 266, 260.2, 257.8, 257.8, 253, 251.4, 241.4, 
    237.4, 237.2, 233, 214.6, 198.8, 200, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  299.7, 293.1, 287.5, 286.9, 285.3, 285.3, 284.7, 281.3, 277.7, 275.3, 
    274.1, 263.6, 262.6, 261.4, 262, 261, 258.2, 252.4, 251.6, 248.2, 241.6, 
    203, 193.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  274.7, 275.1, 265.2, 263.6, 258, 258, 259.2, 258.2, 257.8, 255, 252.4, 
    242.4, 241.4, 239, 238.6, 224.2, 223, 228, 225.2, 227, 223.4, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  282.1, 271, 270.4, 271.4, 272, 272.6, 267.8, 267.4, 266.6, 266.2, 265.6, 
    265.2, 263, 260.8, 256.8, 250.8, 246.6, 233.6, 232.6, 208.6, 214.8, 
    218.2, 220, 220.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  281.1, 282.1, 275.3, 271.4, 268.8, 263.6, 265, 267, 265, 264, 263.2, 262.6, 
    263, 263.6, 263.4, 262.2, 246.4, 245, 239.8, 231.4, 211.4, 219.6, 222.2, 
    220.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  282.5, 278.7, 264.6, 260, 256, 258, 256.2, 255.6, 254.8, 254.6, 254.2, 
    253.2, 252.6, 251, 249.8, 249.6, 246.8, 245.6, 243.8, 236.4, 234.4, 
    226.6, 220.6, 220.2, 224, 222.8, 221.8, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  280.1, 280.7, 283.1, 277.1, 274.7, 274.1, 271.6, 272.8, 273.9, 272.4, 
    270.8, 263.2, 263.6, 255.4, 250.6, 243.8, 230.2, 223.2, 207.8, 216, 
    217.6, 219.6, 220.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  280.5, 280.5, 281.5, 282.1, 274.9, 271.6, 270, 268.4, 254.8, 252.2, 224.2, 
    208.8, 216.2, 219.2, 218.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  283.9, 287.1, 285.9, 287.5, 282.9, 273.1, 258.2, 252.2, 240.8, 234.8, 
    222.4, 208.2, 216, 215.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  297.3, 292.5, 288.5, 289.3, 286.9, 279.9, 276.3, 272.2, 272.4, 267.8, 
    266.8, 264.4, 263.6, 264, 264, 264, 264, 263.4, 262.8, 262, 259.8, 254.4, 
    253.2, 251.6, 250.4, 249.8, 247.4, 246.6, 244.8, 242.6, 238.6, 236.4, 
    233.8, 231.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  292.5, 285.1, 282.9, 275.3, 257.8, 253, 249, 244, 234.6, 231.6, 204, 191.6, 
    194.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  293.5, 295.1, 291.9, 290.3, 290.9, 288.9, 283.7, 283.5, 282.1, 282.3, 
    279.9, 279.9, 279.5, 278.7, 278.5, 276.9, 272.4, 271.8, 268.6, 249, 
    214.2, 206.6, 205.2, 209.6, 209.2, 204.4, 204.4, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  279.9, 273.1, 271.6, 273.7, 269.6, 268.4, 256, 255.2, 252, 249.6, 245.6, 
    243.2, 236.8, 215.2, 212.4, 215, 213.2, 216.8, 214.2, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  283.3, 280.5, 276.7, 278.1, 274.1, 272.8, 270.4, 269, 268.4, 267.6, 266.6, 
    266.4, 266.6, 265.4, 264.6, 263.2, 262.6, 262, 261.8, 261.8, 258.4, 
    258.2, 257.8, 256, 255.8, 249.4, 248.2, 246.2, 224, 213, 217.6, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  300.3, 288.9, 288.1, 287.7, 284.3, 284.5, 280.9, 280.9, 280.1, 278.1, 
    277.1, 273.1, 271.8, 266.2, 265.4, 260.2, 259.8, 258.8, 258.2, 256.2, 
    255, 254.6, 253.2, 249.2, 248.6, 248.6, 245, 244, 240.6, 237.6, 235, 
    212.8, 199.6, 197, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  279.1, 275.1, 275.3, 273.3, 267.4, 268.8, 266.8, 264.8, 260.4, 236.2, 
    224.8, 222, 223.2, 219.2, 220.2, 223.8, 219.8, 221.6, 219.2, 219.6, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  262.4, 264.2, 263, 256.4, 258, 259.2, 259.6, 258.8, 259, 259, 258.4, 257.2, 
    250.8, 247, 244.2, 241, 229.4, 220.6, 220.6, 225.2, 226.2, 228.4, 230.2, 
    229, 231.8, 230, 230.4, 233, 230, 230.8, 228.6, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  295.5, 296.7, 292.1, 290.3, 287.5, 284.7, 282.7, 282.1, 280.9, 281.3, 
    281.5, 279.7, 276.3, 275.9, 275.3, 270.4, 263.2, 215, 204.6, 205.6, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  293.3, 294.3, 292.9, 291.9, 290.7, 290.9, 290.1, 289.9, 288.1, 287.7, 
    281.9, 281.3, 281.7, 279.7, 277.7, 275.5, 266.2, 264.6, 264.6, 264, 
    263.8, 261.2, 260, 255.8, 255.4, 252.8, 251.8, 249.4, 208.2, 201.6, 208, 
    205.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  294.9, 293.7, 294.9, 294.5, 294.3, 293.5, 283.5, 276.1, 273.1, 272.8, 270, 
    269.6, 265.6, 264.6, 263.8, 263, 259.8, 259, 258, 246.2, 240.8, 239, 234, 
    204.2, 202.8, 209.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  294.7, 283.9, 273.1, 272.8, 272.6, 272.4, 269.4, 269, 264.4, 264, 262.4, 
    260.8, 253.4, 252.2, 230, 226.4, 222.2, 206.6, 201, 203.8, 206.4, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  294.9, 294.7, 289.7, 287.1, 281.3, 279.3, 278.5, 278.1, 278.3, 275.7, 
    274.7, 272.4, 271.8, 263.6, 262.4, 259.4, 256.6, 254.4, 251.4, 248.4, 
    247.2, 241.8, 225.4, 202.6, 200.4, 206.4, 208, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  289.1, 283.7, 281.1, 279.1, 275.3, 275.1, 277.1, 275.9, 260.2, 257.6, 
    237.8, 235.2, 206.2, 204.8, 208.4, 203.2, 206.2, 206, 210, 208, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  292.3, 293.5, 278.7, 278.5, 278.5, 273.7, 273.1, 267.6, 267.6, 267, 257.6, 
    242.8, 219.6, 207.4, 201.6, 206.4, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  282.1, 284.3, 285.3, 286.9, 280.7, 280.3, 272, 271.8, 265, 257.8, 247.8, 
    246.6, 233.4, 221.2, 210.6, 207.4, 207.2, 209.6, 211.4, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  288.5, 290.7, 289.9, 284.5, 276.5, 275.9, 275.1, 273.9, 270.6, 271.2, 265, 
    265.2, 263.2, 262.6, 258.4, 239, 213.2, 202, 211.2, 210, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  290.9, 291.3, 291.1, 285.1, 282.9, 280.3, 280.1, 278.5, 274.5, 273.1, 269, 
    263.4, 254.2, 243, 208.2, 205, 205.4, 209, 204.6, 207.8, 210.2, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  279.7, 287.1, 276.1, 274.3, 269, 268.6, 251.6, 251.4, 244.4, 243, 242.4, 
    234.8, 215.4, 211.2, 214, 217.2, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  284.5, 289.1, 276.3, 276.7, 277.1, 266.2, 265.4, 265.2, 264.8, 260.4, 
    261.2, 256.4, 256.4, 247.6, 232.2, 221.6, 216.6, 206.8, 210, 213.6, 212, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  285.3, 288.1, 288.3, 279.1, 280.3, 269, 267.4, 261.8, 219.4, 210, 212.8, 
    210.2, 212.2, 211.2, 214, 217.2, 205.4, 209, 204.6, 207.8, 210.2, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  293.9, 293.5, 295.1, 289.5, 287.3, 282.3, 284.1, 286.1, 271.8, 250, 245.8, 
    226.4, 222.8, 204.4, 199, 205.8, 204, 207.6, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  291.3, 295.5, 293.9, 290.7, 291.1, 290.1, 289.3, 288.7, 282.3, 276.5, 
    276.3, 274.9, 274.7, 268.4, 266, 265.8, 265.4, 264.8, 260.8, 258.2, 
    257.8, 256.6, 254.6, 252.8, 235.6, 210.4, 203, 203, 207.4, 205, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  295.3, 292.3, 292.7, 291.9, 287.3, 285.9, 286.3, 286.5, 273, 267.4, 208.8, 
    202, 203.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  289.5, 290.3, 286.3, 281.5, 281.9, 282.3, 282.9, 286.7, 285.9, 274.9, 
    270.8, 244, 210, 202, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  288.9, 286.7, 291.5, 290.5, 248.2, 239.4, 240.2, 237.2, 216, 204.8, 207.6, 
    202.6, 203.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  292.7, 294.1, 293.5, 290.1, 290.7, 277.9, 275.5, 273.1, 264.6, 261.6, 
    258.6, 259.4, 259, 249.6, 199.8, 207, 205, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  293.5, 294.9, 293.9, 292.7, 293.5, 295.5, 296.5, 294.7, 270.8, 271.4, 
    269.4, 248.6, 233.6, 228.8, 204.4, 201.8, 207.4, 203.6, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  290.5, 292.1, 295.3, 295.7, 292.5, 280.1, 269.4, 266.2, 265, 260.6, 254, 
    250.2, 249, 247.6, 244.6, 236.2, 231.8, 222, 206.2, 205, 209, 205.2, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  297.1, 290.7, 279.3, 265.8, 265.4, 254, 253.6, 251.4, 241.6, 226, 210.4, 
    205.8, 209, 207.4, 202.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  294.5, 287.7, 285.9, 283.1, 273.1, 258.6, 256.8, 257, 258, 256, 251.8, 
    241.8, 235.6, 233.8, 231, 207.4, 212.8, 206.6, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  283.9, 273.1, 272.6, 270.4, 270.2, 268.6, 258.6, 258, 259.4, 245.8, 236.4, 
    234.8, 233, 228, 209.6, 209.4, 216.8, 215.6, 209.4, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  285.5, 278.5, 268.2, 250, 247.6, 245.8, 245.6, 217.2, 220.6, 214.8, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  293.5, 291.9, 292.7, 293.9, 296.7, 287.9, 266.6, 264.2, 263.6, 264, 264.2, 
    257.2, 240.8, 237, 225.8, 213.8, 200, 201, 206, 206.4, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  299.7, 300.1, 273.1, 262.2, 258.2, 255, 251.2, 243.6, 242.4, 239, 237.2, 
    203.6, 209.8, 205.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  278.1, 276.5, 273.3, 271.6, 271.8, 272.8, 272.2, 254.8, 253.8, 254.4, 
    252.2, 246.2, 243.8, 233.4, 208.4, 205.2, 213.6, 210.8, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  293.1, 287.7, 264.6, 263.4, 261.8, 261.6, 261.6, 257, 256.4, 242.4, 209.6, 
    212.6, 210.6, 214.8, 212.8, 212.4, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  282.3, 280.1, 282.5, 280.7, 282.5, 281.7, 281.3, 280.5, 280.1, 278.9, 
    273.1, 273, 271.4, 271.4, 258, 232, 222.6, 220.6, 224.2, 223.8, 216.4, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  293.3, 294.1, 293.5, 289.5, 289.5, 283.7, 278.7, 262.6, 256, 255.6, 242.8, 
    237.2, 234.8, 234.8, 231.2, 224.2, 209.8, 204.2, 210.4, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  283.5, 283.7, 287.5, 287.7, 288.3, 288.9, 285.5, 279.7, 279.1, 277.5, 
    277.9, 255.4, 251.2, 248.6, 249, 248.8, 244, 229.4, 223.2, 220.6, 214, 
    203, 214.6, 210.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  280.9, 282.1, 279.1, 273.1, 268.2, 262, 257.4, 253, 251.8, 251.6, 251.6, 
    234.6, 220.2, 219, 222.2, 216, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  289.1, 290.1, 285.7, 281.9, 274.5, 273, 271.8, 270, 268.4, 267.2, 265.6, 
    265, 264.2, 263.2, 262.8, 251.2, 210.4, 203.8, 212.2, 211.6, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  279.1, 281.1, 279.3, 276.1, 277.1, 276.5, 274.7, 273.9, 273.1, 269.2, 
    267.6, 264.2, 258.8, 251.8, 248, 245.6, 240.4, 233, 233.4, 218, 209.6, 
    214.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  283.5, 283.7, 283.5, 283.3, 282.7, 270.6, 263, 259.2, 253.6, 248.6, 244.4, 
    226.6, 221.2, 220, 222.6, 216.8, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  277.9, 279.3, 275.3, 276.9, 276.7, 270.4, 270.6, 267.2, 264.6, 265.8, 263, 
    258.2, 258, 257.6, 243, 237, 237.4, 236, 224.4, 222.4, 214.2, 220, 218.8, 
    214, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  282.5, 285.7, 287.1, 287.7, 276.3, 266.8, 266.6, 264.4, 264, 259, 247.8, 
    246, 244, 237, 235.2, 232.8, 215.6, 215.4, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  282.9, 283.7, 281.3, 266.8, 263.8, 262.6, 260.8, 258.2, 256.6, 254, 246.4, 
    213.6, 221, 219.2, 217.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  300.1, 294.1, 290.5, 289.9, 288.5, 287.5, 286.5, 286.7, 284.7, 281.7, 
    278.9, 277.1, 277.7, 277.9, 277.5, 277.3, 273.1, 270.2, 269.6, 266.8, 
    260.2, 252.2, 251.4, 251, 216.4, 197, 197.2, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  264, 267, 266.6, 268.6, 264.2, 262.2, 262.8, 259.8, 257.4, 252, 253, 248.8, 
    243.6, 238.4, 233.8, 231, 223.4, 224.2, 222.4, 228, 226.4, 228, 229, 
    230.6, 228.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  280.9, 284.9, 286.9, 284.5, 274.1, 273.1, 271.8, 264.6, 255.4, 245.4, 
    233.4, 224, 214.6, 214, 214.6, 212.4, 215.4, 215.4, 212.4, 215.8, 215, 
    216.6, 215.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  287.1, 279.7, 280.5, 280.5, 269, 259.4, 257.8, 258.6, 254.4, 255, 250.8, 
    247.4, 239.2, 231, 223, 214.6, 211, 211.8, 210.8, 204, 209, 211.2, 213.8, 
    212.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  276.1, 275.1, 278.7, 276.7, 272.4, 268.6, 267.2, 268.2, 269.2, 269.2, 
    265.6, 260.2, 252, 235.2, 222.4, 218.6, 220.6, 223.2, 224, 219.8, 219.2, 
    222.4, 219, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  272.2, 274.5, 273.5, 269.8, 271.4, 264.6, 256.6, 229.4, 214.6, 215.4, 
    220.8, 219.6, 222.8, 225, 224, 225.2, 225.4, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  263.4, 267.4, 269.4, 269.2, 269.4, 269.8, 270, 269, 269.2, 266.6, 252.4, 
    233.6, 222, 219.2, 220.2, 218.8, 222.2, 226.6, 228, 226.2, 227.2, 224.8, 
    226.8, 225, 226.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  291.9, 287.3, 282.1, 278.9, 278.1, 277.9, 278.3, 276.9, 276.9, 276.7, 
    277.3, 273, 261, 259, 253.4, 248.4, 239.6, 236.2, 215.2, 203.6, 203.6, 
    207.4, 204.8, 209.8, 207, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  296.9, 297.1, 293.1, 290.9, 288.1, 282.7, 283.3, 282.1, 273.1, 267, 262.6, 
    262.4, 262.6, 262, 259.8, 258.8, 252.6, 249, 247.4, 245.2, 242.4, 240.2, 
    229, 209, 207.2, 210, 205.4, 205.8, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  294.5, 293.3, 291.9, 292.1, 288.3, 284.9, 283.7, 280.5, 278.7, 272.2, 
    271.2, 254.6, 253, 251.4, 242.8, 236.8, 212.4, 203.4, 206.6, 206, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  295.1, 292.7, 293.9, 290.9, 281.9, 272.6, 269.6, 266.8, 265.2, 256.2, 
    253.4, 241.2, 236.8, 233, 204.6, 201.4, 205.2, 204.6, 208, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  295.1, 289.3, 285.9, 282.7, 277.1, 269.2, 266.6, 266.2, 263.6, 261.4, 
    259.4, 258.8, 252, 242, 208.8, 202.2, 207.6, 205.2, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  292.1, 294.1, 282.5, 276.3, 273.1, 268.4, 266.6, 266.4, 260.8, 254.6, 
    250.2, 249.2, 244.8, 237.2, 225, 213, 201, 201.2, 206.4, 206.4, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  295.9, 291.1, 290.9, 290.9, 290.7, 289.7, 284.3, 283.9, 281.3, 281.3, 
    280.1, 275.3, 274.1, 272, 271.2, 270.6, 268.8, 266.2, 265.2, 262.8, 
    259.4, 253.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  289.9, 289.3, 291.1, 291.1, 289.5, 287.3, 286.7, 284.5, 284.1, 283.1, 
    283.1, 269, 263.6, 259.8, 241.6, 207, 201.6, 200.6, 207, 205, -99999, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  289.9, 291.1, 291.3, 287.3, 275.1, 273.5, 271.6, 272.4, 272.2, 266.4, 
    257.2, 236.2, 233.8, 224.6, 213.4, 200.4, 207.2, 206.2, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  285.7, 287.3, 287.3, 286.7, 286.1, 285.5, 280.3, 280.7, 283.1, 273.7, 
    269.2, 256, 246.6, 245.2, 239.4, 237.4, 215, 207.6, 211.8, 209.4, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  291.1, 283.5, 285.3, 283.9, 282.1, 278.7, 275.9, 273.5, 271.2, 262, 259.2, 
    258.4, 253, 244.8, 213, 209.4, 211.2, 202.8, 209.8, 210.4, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  297.7, 292.1, 289.9, 285.5, 282.7, 281.5, 281.3, 281.9, 277.9, 275.7, 
    273.9, 273.1, 271.4, 270.2, 270.2, 266.8, 263, 262.6, 263, 261.6, 260.8, 
    255, 243.2, 241.6, 235.2, 232, 193.4, 199.4, 208.2, 204.6, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  296.9, 290.5, 288.7, 289.3, 289.1, 284.7, 280.3, 280.3, 279.9, 276.9, 
    270.8, 209, 200.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  296.7, 291.9, 288.3, 288.7, 288.1, 285.7, 283.5, 281.3, 280.9, 280.5, 
    280.1, 278.9, 277.5, 273.1, 256.2, 254, 212.4, 201.6, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  296.5, 289.3, 282.7, 277.9, 277.5, 272, 258.6, 257.6, 236.2, 228.6, 220.2, 
    212.6, 210.8, 207.4, 210, 207.2, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  283.1, 280.9, 280.3, 283.5, 282.5, 282.9, 278.5, 276.7, 273.1, 263.2, 
    263.4, 258, 246.2, 244, 238.4, 236.6, 213.4, 211, 216.6, 217.2, 215, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  276.1, 275.9, 274.7, 269.4, 269, 267.8, 268.2, 249.2, 234.2, 226.4, 221.8, 
    223.4, 217.2, 218.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  287.9, 288.1, 287.1, 282.3, 273.1, 267.4, 265.2, 263.2, 260.2, 258, 257.4, 
    254, 252.8, 250.6, 249.2, 245, 241.8, 237.6, 232.4, 229, 212.6, 211.4, 
    217, 216.4, 215, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  283.7, 281.7, 280.1, 278.9, 277.5, 277.1, 275.7, 269.6, 269, 268.4, 266.2, 
    264.6, 264.2, 263.4, 262.6, 261.6, 261.2, 260.2, 259, 253.4, 238.4, 
    235.6, 229.8, 217.4, 222, 221.4, 216.4, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  284.5, 285.9, 289.1, 289.3, 287.3, 281.5, 274.1, 270.2, 271, 266.2, 265, 
    264.4, 263, 261.4, 256.2, 256.4, 254.8, 254.4, 253.4, 244.8, 244.8, 
    242.2, 203.2, 203.8, 213, 208.6, 212.6, 211.2, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  288.5, 291.1, 282.9, 280.7, 277.7, 277.9, 277.7, 273, 272.4, 273, 270.6, 
    268.8, 264.8, 259, 254.2, 250.8, 250, 246, 233.4, 231.4, 227.6, 225, 
    205.2, 210, 209.2, 213.6, 210.4, 212.4, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  284.7, 278.3, 278.3, 278.3, 280.5, 275.9, 274.5, 270, 267, 258.2, 240.2, 
    221, 207.6, 210.4, 209, 215.2, 212.2, 213.6, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  281.5, 283.3, 281.7, 268.2, 266, 265.4, 263, 258, 256.6, 255.2, 254, 252.8, 
    244.2, 236.4, 233, 228.6, 215.8, 220.6, 217.2, 218, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  279.1, 282.5, 281.7, 281.7, 282.5, 283.5, 260, 259.4, 259.6, 258.4, 257.6, 
    257, 256.6, 252.8, 250.2, 242.4, 233.4, 213.2, 219.4, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  292.1, 288.5, 288.7, 284.3, 285.5, 270.6, 270.8, 268, 244.4, 224.2, 216.6, 
    209.8, 200, 208, 204.4, 205.8, 211.2, 213.2, 219.4, 215.8, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  294.5, 284.3, 284.1, 283.7, 280.7, 279.9, 276.1, 271.6, 269.6, 269.2, 
    263.4, 262.6, 262.2, 262, 261.8, 261.4, 250, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  294.1, 293.9, 292.1, 291.9, 290.9, 290.7, 287.9, 280.3, 279.5, 279.5, 
    279.1, 277.7, 274.3, 274.1, 270.2, 267.8, 266.4, 265.2, 262.8, 262, 
    260.4, 254, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  298.5, 282.5, 281.7, 281.3, 280.3, 279.7, 262.8, 236, 198.6, 190.2, 192, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  262.8, 261.2, 259, 266, 267, 269.8, 269.4, 269.2, 269, 268.4, 267.8, 264.6, 
    252.6, 251.2, 249.2, 239.8, 233.4, 230, 226.2, 217.6, 224.8, 228, 228.6, 
    227, 228.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  279.5, 281.1, 273.9, 274.5, 273.5, 272.2, 271.6, 268, 268.8, 261.2, 255.2, 
    250.4, 248.8, 246.4, 244.6, 241.8, 240.2, 234, 230.4, 212.8, 212.2, 
    215.6, 217.2, 217.6, 219.6, 218.2, 220.2, 219.4, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  278.5, 266.2, 267.2, 268, 268, 263.2, 255.6, 254.6, 249.8, 246.4, 234.2, 
    225.4, 216.8, 216.6, 221, 219.8, 222.8, 222.4, 226.2, 226, 220.8, 221, 
    224.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  265.6, 268.2, 269.4, 271.2, 271.8, 271.4, 271.4, 270.4, 270.2, 269.8, 
    270.8, 268.8, 268, 262.4, 254, 251.8, 234.2, 218.6, 222.4, 225.2, 224.4, 
    219.4, 222.2, 219.6, 220.8, 218.4, 220, 219.6, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  267.4, 263.6, 266.4, 267, 266.8, 257, 255, 254.4, 251.8, 250.8, 249.8, 
    239.8, 227, 219, 220, 222.8, 224, 223, 225.4, 224, 225.6, 224.4, 225.2, 
    222.6, 223.4, 220.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  272.8, 270.4, 267.2, 260.6, 263.4, 263.8, 260.4, 251.8, 250, 246.6, 246.2, 
    241.6, 235, 233.2, 232.4, 226.4, 220.4, 226, 225, 229, 228.6, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  265.8, 266, 262.2, 261.4, 261.6, 264.4, 264.8, 264.2, 262.8, 258.8, 253, 
    248.2, 244.4, 243.8, 241.2, 238.8, 232.4, 226, 221.2, 220.6, 227.4, 
    228.2, 229, 227.2, 228.6, 227, 227.4, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  267.8, 263.2, 264.2, 264.2, 263.8, 263, 262.6, 261.6, 260.2, 259.8, 257.6, 
    255, 253.4, 252.6, 250.2, 248.6, 240.6, 237.6, 234, 220.2, 218.8, 222, 
    220.8, 222.8, 223.4, 225.2, 227.2, 224, 224.6, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  269, 272.8, 272.6, 267, 264.2, 260.4, 259.4, 257, 255.8, 230.8, 220.8, 
    220.6, 222.8, 225.8, 225, 226.4, 229.2, 228, 228.6, 226.2, 227.4, 223.2, 
    224.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  282.9, 270.8, 266.6, 260.2, 259.6, 255.8, 255.2, 255.4, 256, 256.4, 250, 
    249.4, 248.2, 242.4, 239, 236, 230.6, 225.6, 213.2, 216.8, 220.4, 219.4, 
    219.8, 223.4, 219, 221.4, 219.8, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  275.1, 270.6, 271.4, 263.4, 262.2, 245.2, 241.6, 238.6, 224.4, 219.6, 
    223.6, 227.6, 228.8, 225.6, 228.2, 224, 225.8, 223, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  286.7, 271.2, 261.2, 254.8, 252.8, 252.2, 250.4, 242.8, 240.8, 224, 221.4, 
    218.6, 219.6, 217.8, 219.2, 220.6, 216.2, 217, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  299.7, 292.9, 284.1, 281.9, 281.1, 280.5, 278.1, 277.9, 277.3, 274.7, 268, 
    267.8, 266, 263.6, 261.8, 258, 254.4, 239.8, 215.4, 200.2, 196.8, 197.8, 
    197.8, 197.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  284.1, 285.5, 286.3, 279.9, 258, 256.4, 254.8, 253.8, 253.2, 251.2, 244, 
    236.8, 231.8, 229, 225.6, 213.6, 217.6, 220.2, 218.6, 219, 221, 219.4, 
    221, 218.6, 217, 217.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  280.7, 282.9, 279.3, 274.1, 275.1, 273.3, 272.2, 255.8, 235, 227, 225.4, 
    220, 216, 217.4, 213.6, 213.8, 215.4, 216.2, 214.6, 216.6, 215.4, 216, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  264.2, 265.8, 272, 272.6, 268.2, 269.6, 263.8, 263.6, 257.6, 251.6, 237.8, 
    221.4, 219, 221.8, 225.8, 229.2, 225, 226.4, 228, 227.8, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  297.5, 289.3, 289.3, 287.3, 288.7, 290.1, 289.5, 284.9, 279.3, 277.7, 
    273.5, 264.4, 254.2, 233, 207.6, 198.2, 196.4, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  282.5, 278.9, 280.5, 283.1, 285.5, 285.3, 285.7, 273.3, 273, 272.2, 267.6, 
    265.4, 264.8, 263.4, 260.2, 257.6, 248.4, 237, 235.6, 224.4, 208.8, 
    209.4, 216, 217.2, 216, 217, 214.8, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  278.9, 275.7, 270, 269.8, 270.4, 266.8, 263.8, 262, 259.4, 256.8, 254.6, 
    250.6, 249, 231.8, 213.4, 214, 219, 222.4, 221.8, 223.4, 218.6, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  297.5, 297.1, 288.3, 284.7, 285.1, 285.5, 283.3, 283.3, 282.9, 278.5, 
    278.1, 276.1, 275.3, 270, 268.8, 268.6, 263.8, 263.8, 261.6, 258.8, 
    256.4, 255.4, 255.6, 253.4, 245.4, 243.6, 218.6, 214.2, 200, 195.2, 
    195.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  294.3, 289.5, 286.9, 273.1, 271.2, 266.8, 265.4, 264.6, 263.6, 260, 257, 
    252.8, 251.6, 248.6, 246.4, 237, 235.8, 214.4, 213.6, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  297.9, 296.5, 294.5, 293.5, 291.7, 286.3, 285.7, 285.3, 282.5, 281.7, 
    279.9, 279.7, 279.7, 279.5, 277.9, 277.7, 277.5, 277.3, 276.7, 274.9, 
    272.6, 272.6, 272, 270.8, 270, 266.4, 262.6, 261.8, 257.8, 257.2, 255.2, 
    253.8, 253.8, 253.8, 253.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  278.7, 277.3, 276.5, 277.5, 277.3, 277.3, 277.5, 275.5, 269, 269.8, 267.6, 
    263, 259.4, 257.2, 248.8, 237.8, 230.2, 228.6, 222.6, 214.8, 222.6, 
    222.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  285.1, 286.1, 280.5, 281.3, 286.3, 286.7, 283.3, 279.7, 281.1, 281.3, 
    270.6, 261.8, 255.8, 246.6, 231.6, 217.4, 217, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  285.3, 285.1, 286.9, 281.7, 280.5, 263.4, 261.6, 246, 227.6, 216.4, 219.4, 
    216.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  296.5, 297.5, 294.5, 289.3, 285.7, 280.9, 279.7, 277.9, 278.1, 278.5, 263, 
    259, 239, 212.2, 201.4, 201, 196.6, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 tdSigT =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.600006, 3.899994, 4, 3.400024, 6, 8, 17, 17, 21, 21, 18.00002, -99999, 
    -99999, -99999, -99999, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.200012, 2, 0.8999939, 1.5, 4.199997, 3.600006, 5, 29, 29, 28, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.100006, 2, 0.8999939, 1, 0.7000122, 2.5, 2.700012, 3, 9, 32.00002, 
    30.00002, 19, 15, 9, 11, 8, 8, 8, 8, 36.00002, 37.00002, 39.00002, 
    37.99998, 37, 33, 28, 28, 27, 23, 23, 22, 22, 22, 22, 22, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1.5, 3.199982, 1, 1.099976, 1.300018, 2.100006, 6, 8, 15, 28, 19, 11, 6, 6, 
    13, 10, 4, 3.200012, 7, 8, 7, 23, 34, 34, 35, 33, 34, 33, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 2.100006, 7, 3, 5, 3.399994, 0.5, 6, 8, 14, 12.00002, 8, 13, 9, 8, 16, 
    11, 9, 15, 19, 21, 25, 24, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.699982, 0.7999878, 0.8999939, 1, 1, 1.100006, 2.400009, 6, 6, 7, 7, 10, 
    12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.2999878, 0.9000244, 1, 0.3000183, 4.300018, 8, 10, 3, 0.3999939, 
    2.299988, 3, 3, 4, 14, 15, 15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.899994, 0.6000061, 0.7000122, 12, 16, 23, 28, 19, 4.299988, 0.7000122, 
    2.799988, 1.5, 4.300003, 1.899994, 4.800003, 3, 4, 3.600006, 6, 12, 23, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  2.899994, 3.699982, 12, 14, 29, 16, 26, 35.00002, 19, 28, 28, 16, 20.99998, 
    10.00002, 6, 2.600006, 3, 7, 4, 7, 20, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.200012, 3.899994, 1.199982, 4.399994, 1.600006, 7, 11, 9, 20, 13, 32, 26, 
    4.800018, 2.299988, 9, 6.000015, 8.999985, 15.99998, 13, 18, 6, 6, 10, 
    17, 13, 11, 11, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  4.900024, 3.100006, 4.100006, 10, 6, 8, 4.600006, 3.799988, 10, 10, 6, 7, 
    10, 7, 8, 5, 6.000015, 4.5, 9, 10, 3.200012, 4.800003, 5, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1.800018, 1.600006, 0.9000244, 2.800018, 0, 0.6000061, 6.000015, 3.300018, 
    8.999985, 6, 8, 10, 3.299988, 3.800003, 12, 4.099991, 13, 23, 22, 24, 23, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  10, 0.7000122, 1.399994, 17, 12, 15, 10, 21, 13, 19.00002, 16, 30.00002, 
    21, 4.199982, 3.099991, 2, 4.600006, 4.100006, 5, 3.800003, 7, 19, 25, 
    25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  5, 9, 7, 2.100006, 4.299988, 0.8999939, 9, 17, 8, 8, 18.00002, 13, 21, 18, 
    9, 11.00002, 18, 10, 7, 6, 4.099991, 15, 24, 23, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  10, 10, 0.7000122, 0.6000061, 0.8999939, 2, 4.000015, 2.200012, 8, 10, 
    4.699997, 18, 15, 14, 6, 12, 6, 13, 14, 9, 14, 12, 9, 15, 21, 23, 23, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.200012, 3.400024, 6, 4, 0.7000122, 6, 10, 18.99998, 14, 6, 8, 1.800018, 
    3.800018, 2.799988, 4.400009, 4.900009, 1.699997, 2.800003, 3.600006, 7, 
    15, 22, 22, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  2.5, 0, 15, 17, 31, 13, 16, 11, 4.600006, 7, 3, 3.100006, 10, 23, 23, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.699982, 6, 7, 9, 8, 19, 7.000015, 8, 8, 4.100006, 5, 5, 6, 8, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  4.599976, 0.7999878, 1.100006, 6, 6, 4.799988, 1.299988, 0.8000183, 
    3.799988, 0.5999756, 0.6999817, 7, 18, 8, 14, 40, 9, 19, 16.99998, 7, 
    11.99998, 10, 6, 10, 7, 11, 2.799988, 10, 10, 4.300003, 2.600006, 7, 5, 
    11, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.399994, 2.800018, 8, 7, 0.7999878, 1.399994, 5, 3.399994, 6, 11, 
    4.399994, 3.900009, 4.100006, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.5, 3.600006, 7, 4.799988, 11, 4.199982, 4.400024, 12, 14, 23, 19, 30, 18, 
    16, 28, 34, 18, 23.99998, 20, 25, 8, 8, 8, 9, 10, 12, 12, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 0.3000183, 0.3000183, 4.100006, 2.800018, 4.799988, 2.100006, 4.099991, 
    3, 10, 6, 1, 3.600006, 2.599991, 4.399994, 5, 16, 18, 19, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  3.399994, 0.8999939, 0.9000244, 7, 8, 25.99998, 21, 9, 11, 8, 8, 23, 12, 
    13, 39, 11.00002, 24, 15, 37.99998, 39.99998, 39, 12.00002, 6.999985, 16, 
    38, 32, 10, 9, 8, 8, 13, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  2.5, 5, 2.200012, 4.700012, 2.299988, 8, 3.899994, 8, 8, 3.200012, 9, 7, 
    12, 6, 12, 8.000015, 16.99998, 19.99998, 4.600006, 1.800018, 1.899994, 6, 
    8, 0.3999939, 0.4000092, 3.300003, 4.300003, 16, 18, 13, 3.399994, 
    3.600006, 4.400009, 4.600006, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  3, 3.600006, 4.899994, 8, 3.899994, 12, 26.99998, 32.99998, 34, 20, 14, 13, 
    19, 20, 24, 27, 29, 33, 33, 33, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 1.900024, 2.799988, 0.5999908, 7, 9.000015, 6, 3.599991, 7, 4.600006, 
    2.699997, 5.000015, 5, 19, 15, 6, 4.399994, 4.100006, 8, 16, 23, 25, 31, 
    31, 37, 36, 36, 37, 36, 36, 36, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  3.799988, 5, 1.700012, 7, 7, 17, 15, 7, 7, 19, 21, 34.00002, 32.99998, 15, 
    31.99998, 17, 23.00002, 13, 15, 15, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5999756, 1.299988, 1.5, 13, 7, 14, 10, 17, 7, 12, 6, 7, 14, 10, 25.00002, 
    27, 3.300018, 2.800018, 10, 14, 38.99998, 32.00002, 10, 10, 17, 17, 36, 
    36, 10, 9, 10, 10, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.799988, 3.700012, 10, 10, 3.699982, 6, 1.299988, 6, 3.700012, 8, 
    3.600006, 6, 4.200012, 7, 4.099976, 7, 5.999985, 17, 28, 19, 6, 16, 17, 
    4.5, 6, 12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  7, 3.799988, 4.100006, 4.799988, 12, 7, 7, 12, 7, 11, 11, 20.99998, 19, 25, 
    12, 6, 9, 5, 4.899994, 5, 11, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.799988, 2.800018, 1.300018, 8, 8, 5, 0.7999878, 1.399994, 10, 13, 
    2.900024, 3.100006, 7, 17, 3.600006, 14, 7, 8, 15, 10, 15, 8, 4.299988, 
    6, 6, 6, 7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.6000061, 4.700012, 2.200012, 7, 7, 8, 47, 44, 41.00002, 40, 23, 6, 
    4.599991, 4.5, 4.899994, 5, 5, 5, 6, 12, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.2999878, 1.899994, 3.900024, 2.299988, 5, 10, 18, 14, 10, 13, 8, 14, 5, 
    4.599991, 4.600006, 9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.6000061, 1.799988, 5, 8, 7, 15, 15, 15, 12, 12.99998, 4.600006, 4.800003, 
    4.799988, 3.899994, 3.5, 3.199997, 3.199997, 3.600006, 23, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.7999878, 0.8000183, 4.600006, 0.7999878, 1.600006, 5, 10, 12, 4.899994, 
    14, 17, 32.00002, 37.00002, 33, 14, 15, 8, 7, 8, 8, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 1.199982, 2.899994, 0.5, 4.799988, 8, 13, 11, 7, 13, 8, 3, 1.300003, 
    2.600006, 3.199997, 3.399994, 3.5, 3.899994, 4.300003, 4.900009, 7, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  4.100006, 13, 9, 16, 20, 15, 19, 21, 11, 4.5, 4.299988, 4.699997, 6, 6, 6, 
    8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 16, 10, 15, 22, 22.00002, 36, 18.00002, 28.99998, 24, 33.00002, 27, 11, 
    9, 11, 8, 9, 4.800003, 6, 18, 19, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.099976, 14, 14, 13, 27.99998, 30, 39, 28.99998, 11, 7, 7, 10, 17, 6, 6, 
    8, 3.5, 3.899994, 4.300003, 4.900009, 7, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.399994, 2.200012, 3.800018, 1.200012, 5, 1.599976, 16, 26, 34.99998, 19, 
    23, 12, 6, 4.799988, 4.800003, 6, 8, 10, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.199982, 0, 5, 6, 13, 17, 11, 12, 11, 6, 11, 9, 13, 13, 11, 18.99998, 17, 
    7, 4.799988, 6.000015, 10.99998, 7, 18, 13, 19, 11, 9, 9, 10, 15, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.399994, 0.7999878, 8, 9, 10, 6, 10, 23, 20, 35, 9, 9, 12, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.7000122, 0.6999817, 0.6999817, 6, 5, 31.99998, -99999, -99999, -99999, 
    -99999, -99999, 34, 11, 10, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.299988, 2, 27, 44, 26, 11, 14, 22, 6, 10, 11, 12, 13, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0, 2.200012, 7, 5, 24, 8, 13, 10, 4.800018, 7, 8, 12, 13, 15, -99999, 
    -99999, -99999, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.100006, 4.299988, 7, 5, 7, 26, 31, 30, 13, 21, 31, 26, 8, 15, 6, 5, 9, 
    11, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.799988, 11, 35, 35, 29, 17, 4.5, 14.00002, 11, 19, 19, 22, 11, 20, 21, 
    19, 7, 10, 4.800003, 5, 9, 11, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  16, 24, 17, 4, 11, 18, 33, 27, 13, 11, 11, 11, 12, 14, 14, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  20, 16, 25, 16, 13, 2.399994, 4.999985, 12, 14, 14, 13, 11, 9, 4.800003, 9, 
    7, 7, 7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  18, 6, 8, 6, 25.00002, 24, 3.300003, 4.399994, 16, 6, 8, 2.800003, 
    1.300003, 3, 2.700012, 3, 6, 13, 14, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  19, 18, 26.00002, 15, 3.5, 6, 12, 8, 9, 9, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  2.200012, 4.899994, 10, 17, 25, 19, 1.5, 2.100006, 6, 13, 16.00002, 
    31.00002, 20, 8, 10, 5, 6, 6, 8, 11, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  16, 17, 9, 2.700012, 2.600006, 16, 15, 8, 3.699997, 3.100006, 6, 5, 6, 6, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6, 0.6000061, 0.09997559, 0.3000183, 0.2999878, 9, 12, 2.199997, 4.699997, 
    12, 26, 22, 8, 3.099991, 3.599991, 4.599991, 8, 14, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  25, 18, 1.700012, 3.799988, 18.99998, 20, 7, 5, 1.299988, 7, 6, 7, 13, 16, 
    18, 18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.7999878, 0.8000183, 5, 12, 7, 10, 17, 25, 14, 22, 17, 43, 26, 42, 38, 27, 
    22, 20, 25, 27, 25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.5, 9, 17, 11, 18, 13, 20, 2.800018, 4.600006, 9, 14, 12, 7, 4.900009, 8, 
    5, 6, 7, 14, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 6, 14, 11, 5, 14, 16, 11, 6, 5, 18, 7, 1.300003, 3.400009, 15, 22, 24, 
    10, 16, 9, 4.300003, 4, 12, 15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  9, 8, 10, 7, 1.900024, 1.299988, 4.099991, 3, 6, 14, 16, 12, 10, 10, 11, 
    10, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1.200012, 1.600006, 11, 8, 3.899994, 0.7999878, 0.7000122, 13, 17.00002, 
    12, 17, 12.00002, 23.00002, 16.99998, 29, 11, 9, 11, 12, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.5, 3.600006, 3.899994, 6, 13, 15, 15, 27, 20, 18.00002, 37, 36.00002, 
    12.99998, 8, 1.699997, 1.300003, 9, 8, 13, 8, 8, 19, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  9, 6, 2.799988, 10, 7, 14, 17, 12.00002, 31, 35, 15, 16, 27, -99999, 
    -99999, -99999, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 2.199982, 2.399994, 7, 8, 8, 15, 10, 12, 26.99998, 23, 15.00002, 26, 24, 
    17, 10, 19, 23, 9, 10, 16, 21, 23, 22, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.700012, 7, 7, 11, 10, 4.899994, 9, 3, 10, 16, 11, 3.600006, 2, 2.899994, 
    9, 11, 8, 8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.699982, 6, 7, 0.6999817, 1.799988, 6, 3.799988, 14.00002, 14, 6, 13, 8, 
    15, 26, 25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 5, 3.200012, 0.7999878, 3.600006, 1.100006, 6, 11, 11, 5, 10, 6, 
    29.00002, 40, 30, 16, 18, 11, 17, 9, 17.00002, 7, 14, 11, 11, 7, 7, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.799988, 1.200012, 0.3000183, 3.899994, 1.600006, 3.200012, 2, 1.199982, 
    3.899994, 2.5, 6, 6, 8, 5, 9, 7, 11, 13, 15, 26, 28, 28, 31, 32, 31, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.8999939, 8, 13, 15, 7, 18, 13, 30, 23, 28, 11, 11, 9, 9, 10, 11, 14, 17, 
    19, 22, 23, 24, 25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  11, 12, 24, 23, 32, 27, 2.999985, 1.700012, 1.099991, 6, 10, 8, 9, 5, 6, 6, 
    7, 7, 8, 8, 9, 10, 16, 19, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.8999939, 1.300018, 4.800018, 9, 11, 5, 8, 15.00002, 28.00002, 26.00002, 
    18, 22.00002, 25, 14, 10, 11, 18, 22, 30, 29, 29, 29, 28, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.600006, 8, 10, 5, 0.6999817, 1.899994, 2.800003, 4, 3.800003, 4.799988, 
    10, 16, 20, 27, 27, 27, 27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.1000061, 0, 0, 2.300018, 22, 28.99998, 15, 1.5, 1.400024, 2.300018, 2, 
    2.800003, 6, 7, 8, 9, 11, 17, 18, 18, 19, 18, 19, 20, 22, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.199982, 0, 0.5, 0.1999817, 3.300018, 4, 10, 7, 14, 13, 25.99998, 28, 11, 
    24, 12, 6, 9, 6, 6, 5, 5, 6, 7, 9, 10, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.199982, 4.399994, 1.700012, 2.299988, 14, 12, 29.99998, 36, 29, 25, 10, 
    10, 21, 20, 11.99998, 15.99998, 8, 15, 12, 18, 17, 10, 10, 8, 8, 9, 8, 8, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.399994, 8, 7, 13, 1.799988, 1, 6, 3, 7, 12, 21.00002, 22, 13, 20, 9, 12, 
    7, 6, 7, 12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.3999939, 0.7000122, 12, 1.100006, 4, 3.600006, 5, 8, 9, 6.000015, 11, 11, 
    9, 17, 11, 11, 12, 15, 18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.800018, 6, 3.299988, 6, 2.5, 4.5, 4, 7, 4.300018, 7, 4.299988, 6.999985, 
    10, 16, 9, 7, 10, 12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 3, 3.399994, 4.699982, 16, 13, 16, 10, 19.99998, 14, 25, 13, 21, 9, 12, 
    8, 7, 7, 9, 13, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.600006, 2.200012, 15, 12, 18, 11, 11, 25, 18, 30.99998, 15, 8, 25, 18, 6, 
    13, 8, 10, 20.00002, 14.99998, 31, 22, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0.8000183, 5, 9, 7, 12, 10, 6, 8, 23, 20, 32, 10.99998, 18, 8, 7, 7, 
    10, 10, -99999, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 3.100006, 4.599976, 2.5, 4.700012, 9, 5, 20, 21.00002, 14, 25.00002, 10, 
    4.100006, 11, 6, 4.599991, 8, 10, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 12, 15, 4.900024, 4.700012, 13, 10, 22, 40, 34.00002, 40.00002, 24, 
    21, 13, 10, 3.699997, 3.300003, 6, 13, 17, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.600006, 1.100006, 17, 8, 20, 18, 40, 41, 14, 15, 11.00002, 5, 10, 4.5, 
    4.600006, 5, 6, 7, 10, 15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.200012, 0.8000183, 2.600006, 0.7999878, 0.8000183, 1.5, 4.5, 8, 1.100006, 
    3.900024, 0.8999939, 6, 7, 2.700012, 5, 0.7999878, 1.100006, 3.600006, 
    11, 19, 13.99998, 14, 5, 16, 8, 11, 6, 7, -99999, -99999, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.399994, 1.5, 4.400024, 17, 15, 9, 12, 30.99998, 46, 45, 37.99998, 12, 10, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.400024, 1.5, 6, 15, 13, 9, 13, 9, 32, 33, 19, 15, 45, 41, 25.00002, 30, 
    12, 10, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  24, 31, 30.00002, 17, 28, 27, 15, 29, 12, 4.900009, 7, 6, 12, 13, 16, 16, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.7000122, 0.8999939, 11, 16, 46, 47, 45, 13, 15, 11.00002, 40, 38, 11, 17, 
    11, 24, 13, 13, 15, 17, 16, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.700012, 0.1999817, 5, 1.399994, 6, 7, 16.00002, 24, 7, 9, 18, 26, 24, 24, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  12, 13, 16, 20, 16, 8, 4.300018, 6, 2.900024, 6, 3.299988, 2, 10, 10, 4, 
    3.300003, 8, 2.800003, 3.399994, 12, 8, 7, 15, 22, 22, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.400024, 6, 1.399994, 2.299988, 11, 8, 4.300018, 4, 6, 3.600006, 3.700012, 
    5, 2.700012, 9, 12, 2.399994, 1.900024, 4.500015, 1.799988, 3.5, 5, 8, 
    4.5, 4.899994, 9, 27, 25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.6000061, 0, 0, 0, 4.699982, 1.700012, 0.7000122, 2.300018, 5, 0, 
    1.899994, 4.600006, 7, 2.299988, 2.900009, 8, 6, 12, 14, 7, 4.199997, 
    2.599991, 3.599991, 3.699997, 5, 7, 9, 12, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 12, 14, 8, 11, 22, 20, 13, 17, 37, 14, 12.99998, 7, 11, 5, 8, 5, 14, 13, 
    18, 7, 5, 5, 7, 9, 11, 16, 18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  7, 2.5, 8, 11, 18, 11, 10, 3.799988, 6, 1, 2.800003, 8, 8, 9, 10, 12, 14, 
    18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 6, 7, 1.600006, 8, 3.799988, 6, 9, 4.400009, 3.899994, 11, 9, 10, 4.5, 
    9, 8, 10, 14, 20, 12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2.5, 4.200012, 2.900024, 14, 17, 6, 7, 39, 29, 13, 12, 19, 37, 22, 33, 
    11, 8, 10, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.5, 0.7999878, 4.400024, 4, 16, 15, 30.99998, 35, 24, 10, 11, 6, 5, 7, 9, 
    11, 13, 8, 10, 12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5, 2.799988, 0.7000122, 3.300018, 4.800018, 2.199982, 4, 4.5, 1.700012, 
    4.600006, 3.699982, 14, 9.000015, 14, 9.999985, 39, 36, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  6, 12, 9, 14, 8, 15, 4.5, 7, 3, 8, 5, 10, 3.699982, 8, 6, 11, 8, 11.00002, 
    7.999985, 12, 6, 12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.200012, 4.100006, 9, 6, 10, 11, 29.99998, 30, -99999, -99999, -99999, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.8999939, 0.1000061, 0, 3.399994, 10, 15.99998, 23, 16.00002, 13, 18, 10, 
    5, 7, 12, 9, 14, 7, 9, 5, 3.900009, 12, 31, 36, 35, 36, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8, 12, 10, 11, 13, 9, 3.5, 1.200012, 4.099976, 7.000015, 4.5, 6, 10, 8, 17, 
    13, 5, 4, 6, 4.900009, 6, 9, 17, 22, 24, 26, 26, 29, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  10, 3.400024, 8, 9, 16, 12.00002, 26, 18, 11, 15, 4.199997, 9, 8, 8, 10, 
    13, 17, 23, 35, 35, 33, 33, 34, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.8000183, 5, 2.299988, 0, 0, 0, 3.799988, 9, 11, 21.99998, 26.99998, 
    25.99998, 15, 19, 17, 15, 15, 11, 15, 24, 25, 26, 27, 26, 26, 26, 26, 26, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8, 6, 11, 13, 12.99998, 22, 21, 10, 7, 15, 10, 14, 7, 7, 10, 12, 13, 14, 
    17, 18, 20, 20, 23, 23, 25, 24, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.599976, 2.600006, 4.100006, 0, 1.600006, 3.399994, 10, 10, 20, 19, 19, 
    16, 3.899994, 5, 8, 10, 9, 19, 23, 31, 31, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.299988, 4.200012, 0.6000061, 0.1000061, 0, 0, 8, 6, 4.299988, 8.999985, 
    3.300003, 9, 6, 13, 16, 8, 13, 10, 9, 10, 23, 28, 28, 31, 31, 31, 31, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  7, 9.000015, 15.00002, 12.00002, 17.99998, 12, 18, 12, 20.00002, 15.99998, 
    21, 20, 9, 18, 19, 7, 10, 8, 13, 6, 5, 9, 11, 12, 17, 20, 28, 27, 27, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 6, 6, 1.600006, 8, 6, 9, 2.5, 2.199997, 4.300003, 7, 10, 12, 16, 
    18, 19, 19, 18, 19, 18, 18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  11, 3.799988, 0, 0.4000244, 2.600006, 0.5, 2.699997, 11, 20, 14, 15, 29, 
    26, 22, 5, 2.600006, 5, 4.400009, 2.699997, 10, 18, 23, 26, 30, 29, 31, 
    31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.200012, 0.3000183, 2.5, 0.1000061, 2.800018, 2.800003, 12, 15, 4.299988, 
    4.700012, 12, 24, 31, 30, 35, 34, 35, 34, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  9, 0.4000244, 1, 4.5, 4.699997, 1.899994, 3.5, 3.199997, 5, 2.800003, 
    3.099991, 8, 9, 11, 11, 11, 11, 9, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.700012, 2.5, 47, 35, 1.100006, 0.8999939, 17, 0.5, 0.5, 49.00002, 28, 
    3.699982, 2.299988, 9, 5.999985, 2.5, 18, 6, -99999, -99999, -99999, 
    -99999, -99999, -99999, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.100006, 6, 8, 7, 0.1000061, 1.299988, 7, 6, 16, 17, 3.899994, 8, 8, 10, 
    4.100006, 2.600006, 9, 12, 17, 19, 21, 21, 23, 22, 24, 24, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.600006, 12, 17, 13, 20, 39.99998, 28.00002, 25, 21, 19, 11, 5, 6, 8, 12, 
    13, 14, 19, 19, 24, 25, 28, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 6, 12, 14, 13.00002, 16, 13.99998, 21, 19, 21, 14, 11, 11, 16, 22, 36, 
    34, 35, 35, 35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  3.299988, 9, 14, 10, 27, 36, 38, 19, 14, 24.00002, 21, 21, 2, 32, -99999, 
    -99999, -99999, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.100006, 0, 0, 7, 13, 14, 21, 13, 22, 14, 13, 29, 13.99998, 11, 10.00002, 
    7, 11, 5, 8, 4.5, 4.100006, 4.099991, 9, 16, 21, 28, 31, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  9, 4.5, 0.3999939, 1.299988, 2.5, 2.099976, 11.99998, 10, 25, 16.99998, 8, 
    7, 3.199997, 3.100006, 4, 4.899994, 12, 25, 27, 27, 26, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1, 1.100006, 1.099976, 4.400024, 7, 4.399994, 1.099976, 3.099976, 3.399994, 
    7, 13, 10, 6, 3.200012, 2.099976, 0.3999939, 1.299988, 1.899994, 6, 
    3.399994, 10, 9, 6, 4.599991, 6, 7, 11, 13, 10, 9, 9, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  29, 19, 16, 15, 16.00002, 9, 7, 13, 10, 11, 17, 23, 12, 7, 4.399994, 6, 7, 
    -99999, -99999, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6, 7, 6, 6, 8, 6, 3.900024, 10, 4.100006, 8, 4.299988, 7, 3.5, 2.899994, 
    4.5, 10, 7, 10, 11, 6, 8, 12, 6, 11, 9, 45, 12, 11.99998, 8.999985, 
    8.000015, 12, 3.199997, 3.199997, 3.199997, 3.199997, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.800018, 6, 2.299988, 7, 9, 5, 9, 3.600006, 1.200012, 2.5, 4.200012, 2, 7, 
    3.700012, 8, 11, -99999, -99999, -99999, -99999, -99999, -99999, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  4.300018, 4.300018, 1.100006, 4.399994, 15, 18, 11, 9, 30, 27.99998, 31, 
    45.99998, 39, 24, -99999, -99999, -99999, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  7, 7, 12, 12, 32, 31, 31, 26, 19, 17, 18, 17, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1.600006, 1.899994, 2.600006, 4.799988, 1.100006, 3.399994, 9, 3.199982, 
    37, 37, 32, 33, 28, -99999, -99999, -99999, -99999, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _ ;

 htSigW =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 1500, 1800, 2100, 2400, 2700, 3000, 3300, 3600, 3900, 4200, 4500, 4800, 
    5100, 5400, 5700, 6000, 6600, 7200, 7800, 8400, 9000, 9600, 10200, 10500, 
    11400, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 
    5100, 6000, 7500, 7800, 9000, 10500, 11100, 13200, 15000, 15900, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 
    6000, 7200, 7500, 8400, 9000, 10200, 10500, 11100, 11400, 12300, 13200, 
    13500, 13800, 14100, 14400, 15000, 15300, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    6300, 7500, 8400, 9000, 9600, 10500, 11400, 12000, 12300, 12900, 14700, 
    15000, 16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 
    5400, 6000, 7500, 9000, 9600, 10500, 14100, 15000, 15900, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 9300, 10500, 10800, 15000, 15900, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 7200, 7500, 
    9000, 9900, 10500, 11400, 13200, 15000, 15900, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5100, 
    6000, 6300, 7500, 9000, 9300, 10500, 12000, 13500, 15000, 16200, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 10500, 11400, 12600, 14400, 15000, 15900, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 8700, 9000, 10500, 10800, 12000, 14700, 15000, 16200, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 
    4800, 5700, 6000, 6300, 6900, 7500, 7800, 9000, 9600, 10500, 12300, 
    13200, 15000, 16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 10500, 10800, 11100, 13200, 14400, 15000, 15300, 16500, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 8700, 9000, 10500, 11400, 12300, 15000, 15900, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 10500, 11700, 12900, 15000, 15900, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 
    6000, 7500, 9000, 10500, 10800, 12600, 15000, 15900, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4800, 
    6000, 7500, 9000, 10500, 11700, 12900, 15000, 15300, 15900, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 
    5400, 6000, 7500, 8100, 9000, 10500, 12000, 12900, 15000, 16200, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 4800, 
    6000, 7500, 9000, 10500, 11100, 14700, 15000, 15600, 15900, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3000, 3600, 3900, 4200, 
    4800, 5400, 6000, 7500, 9000, 10500, 12000, 14700, 15000, 15900, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 
    6000, 7500, 7800, 9000, 10500, 11700, 12600, 13500, 15000, 15300, 16200, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4800, 
    5700, 6000, 7500, 7800, 9000, 10200, 10500, 10800, 11100, 11700, 12900, 
    15000, 15600, 16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 4800, 
    6000, 7500, 9000, 10500, 11700, 12300, 13500, 15000, 15900, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 1800, 2100, 2400, 2700, 3600, 4200, 4500, 4800, 6000, 7500, 9000, 10500, 
    11400, 14400, 15000, 15600, 16200, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 
    6000, 6300, 7500, 8400, 9000, 10500, 11100, 12300, 13500, 15000, 15900, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4800, 
    5700, 6000, 6600, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 
    4800, 6000, 7500, 9000, 10500, 12600, 12900, 13800, 14400, 15000, 15300, 
    15600, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4500, 4800, 
    6000, 6900, 7500, 9000, 9300, 10500, 10800, 11700, 12300, 12600, 13200, 
    15000, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4500, 
    4800, 6000, 7500, 9000, 9900, 10500, 12000, 12900, 13500, 15000, 15900, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4800, 
    5400, 6000, 6300, 7200, 7500, 7800, 9000, 10200, 10500, 11400, 12900, 
    13500, 14100, 14700, 15000, 15300, 16200, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3000, 3300, 3600, 4200, 
    4800, 6000, 7500, 7800, 8700, 9000, 10500, 13500, 14700, 15000, 16200, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 6000, 7500, 
    9000, 10200, 10500, 10800, 12600, 13800, 15000, 15300, 16200, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 
    4800, 5700, 6000, 7200, 7500, 8100, 8700, 9000, 10200, 10500, 13200, 
    14100, 15000, 15300, 16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4500, 4800, 
    6000, 7500, 9000, 9600, 10500, 11700, 13200, 14100, 14400, 15000, 15600, 
    16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 600, 900, 1200, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 4500, 4800, 
    5100, 6000, 7500, 9000, 9600, 10500, 11400, 13500, 15000, 15300, 15900, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 
    4800, 6000, 6900, 7500, 9000, 10200, 10500, 11400, 12300, 12600, 13200, 
    13500, 15000, 15300, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 4800, 
    5400, 6000, 7500, 8700, 9000, 10500, 12300, 13800, 15000, 15300, 15900, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4500, 
    4800, 5400, 6000, 6300, 7500, 9000, 10500, 11100, 12600, 13500, 14400, 
    15000, 15300, 16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5700, 6000, 7500, 
    9000, 10500, 10800, 12300, 13200, 15000, 15900, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5400, 
    6000, 6900, 7500, 9000, 10500, 11700, 12600, 12900, 15000, 15300, 15900, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 7800, 9000, 10500, 10800, 12900, 13800, 15000, 15900, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4800, 
    6000, 7500, 8400, 9000, 10500, 11700, 12300, 13800, 14100, 14400, 14700, 
    15000, 15300, 16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 9900, 10500, 12300, 12900, 13500, 14400, 15000, 16200, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 7500, 9000, 
    9600, 10500, 11400, 12900, 14100, 14700, 15000, 16200, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5100, 5700, 6000, 
    6300, 6900, 7500, 8400, 9000, 10500, 11400, 12900, 15000, 15900, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 9900, 10500, 13200, 13800, 14700, 15000, 16200, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 4200, 4500, 4800, 
    6000, 7500, 8100, 8400, 9000, 9300, 10500, 11100, 12000, 14400, 15000, 
    15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 1200, 1500, 1800, 2100, 2400, 2700, 3000, 3300, 3600, 4200, 4800, 5400, 
    6000, 7500, 9000, 10500, 10800, 12000, 14100, 15000, 15900, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 1800, 2100, 2400, 2700, 3600, 4200, 4500, 4800, 5100, 6000, 6900, 7500, 
    8700, 9000, 10200, 10500, 11100, 12600, 13200, 13500, 14700, 15000, 
    16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4800, 5400, 6000, 7200, 7500, 
    8100, 9000, 9600, 10500, 11400, 12900, 13800, 14700, 15000, 16200, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 2400, 2700, 3600, 4200, 4800, 6000, 7500, 9000, 9600, 10500, 12300, 
    14400, 15000, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 3900, 4200, 4800, 6000, 7500, 
    9000, 10200, 10500, 12300, 12900, 13500, 14700, 15000, 15900, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 
    5400, 6000, 7500, 9000, 9300, 10500, 11400, 12900, 13800, 14700, 15000, 
    16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 6900, 
    7500, 8100, 9000, 9900, 10500, 13500, 15000, 15300, 15900, 16200, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 6900, 7500, 9000, 10500, 
    12000, 15000, 16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 6000, 7500, 8400, 9000, 
    10500, 11100, 11700, 14700, 15000, 16200, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4800, 
    6000, 6600, 7500, 9000, 9300, 10500, 11700, 13200, 15000, 16200, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4500, 4800, 6000, 
    6300, 7500, 8400, 9000, 9900, 10500, 12300, 13500, 15000, 15300, 15900, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 3900, 4200, 4800, 6000, 
    7500, 7800, 9000, 10500, 12600, 13500, 15000, 15900, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 2400, 2700, 3600, 4200, 4800, 6000, 7500, 9000, 10500, 10800, 12900, 
    13800, 15000, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 
    5400, 6000, 7500, 9000, 10500, 12600, 13800, 15000, 15900, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 600, 900, 1200, 1800, 2100, 2400, 2700, 3000, 3300, 3600, 3900, 4200, 
    4800, 5100, 6000, 7500, 7800, 9000, 10500, 12000, 13500, 15000, 15900, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 5400, 6000, 
    7500, 8100, 9000, 9900, 10500, 12000, 15000, 15900, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4500, 4800, 6000, 
    7500, 7800, 9000, 9600, 9900, 10500, 11400, 13200, 13500, 15000, 15900, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 900, 1200, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4800, 6000, 6300, 
    7500, 9000, 9300, 10500, 11100, 13200, 14700, 15000, 15900, 11400, 12300, 
    15000, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5700, 6000, 7500, 
    7800, 8700, 9000, 9600, 10500, 12900, 13800, 15000, 15900, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5700, 
    6000, 7500, 9000, 9600, 9900, 10500, 10800, 12600, 13500, 14400, 15000, 
    16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 
    6000, 6900, 7500, 8100, 9000, 10200, 10500, 11100, 12000, 12300, 12600, 
    12900, 13200, 13500, 13800, 14100, 14400, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 
    4800, 6000, 6300, 7500, 9000, 10200, 10500, 14400, 15000, 15900, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 
    6000, 6600, 7500, 8400, 9000, 10500, 11700, 13200, 14400, 15000, 15600, 
    16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3000, 3300, 3600, 
    4200, 4800, 6000, 7500, 9000, 9600, 10200, 10500, 11700, 13200, 13800, 
    14700, 15000, 15300, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5100, 
    5700, 6000, 6600, 7500, 8100, 9000, 9900, 10500, 12300, 13800, 15000, 
    15300, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4500, 
    4800, 6000, 6900, 7500, 9000, 9900, 10500, 11100, 11700, 14100, 14400, 
    15000, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 4800, 
    6000, 6600, 7500, 9000, 9300, 10500, 10800, 12000, 15000, 15900, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 10500, 13200, 14400, 15000, 16200, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 8400, 9000, 10500, 11100, 11700, 12300, 13200, 13500, 14100, 15000, 
    16200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3000, 3300, 3600, 
    3900, 4200, 4500, 4800, 5100, 5400, 5700, 6000, 6300, 6900, 7500, 8100, 
    8400, 9000, 10200, 10500, 13500, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 4200, 4800, 6000, 7500, 9000, 9600, 10500, 10800, 
    12300, 15000, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4800, 
    6000, 7500, 9000, 9300, 10500, 11700, 13500, 14100, 14400, 15000, 15900, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 
    5700, 6000, 6600, 7200, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 3900, 4200, 
    4800, 5100, 6000, 7200, 7500, 7800, 9000, 10500, 12000, 14100, 14400, 
    15000, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4500, 4800, 
    5400, 6000, 6900, 7500, 8100, 8700, 9000, 9600, 10200, 10500, 12000, 
    12900, 15000, 15300, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 
    4500, 4800, 6000, 7500, 8400, 9000, 10500, 11100, 13200, 14700, 15000, 
    15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 7500, 
    8400, 9000, 10500, 12300, 13500, 13800, 15000, 15900, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5400, 
    5700, 6000, 7500, 8700, 9000, 9900, 10500, 10800, 12000, 12900, 14400, 
    15000, 16200, 14100, 14400, 14700, 15000, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 9600, 10500, 12600, 15000, 15900, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    6600, 7500, 8100, 9000, 9300, 10500, 11700, 13800, 15000, 16200, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5700, 6000, 7500, 
    9000, 9300, 10500, 12000, 12300, 13200, 13800, 15000, 15900, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 9900, 10500, 11400, 14100, 15000, 15900, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 6000, 6600, 7500, 9000, 
    10500, 11100, 12000, 14400, 15000, 15900, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 1500, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 7500, 9000, 10500, 
    11100, 12600, 13500, 15000, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5400, 6000, 
    7500, 9000, 9600, 10500, 10800, 15000, 15900, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4800, 
    5100, 5700, 6000, 7500, 9000, 9300, 10500, 12000, 13800, 15000, 15900, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 
    6000, 7500, 8700, 9000, 10500, 12000, 13500, 14700, 15000, 15300, 15900, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 7500, 9000, 10500, 
    11700, 15000, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 1200, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 4800, 5100, 6000, 7500, 
    7800, 9000, 9900, 10500, 12000, 12900, 14100, 15000, 15900, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 
    4800, 5100, 5700, 6000, 7500, 9000, 9600, 10500, 11100, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3000, 3600, 3900, 4200, 
    4800, 6000, 7500, 9000, 10500, 12600, 13200, 15000, 15900, 12600, 12900, 
    13200, 15000, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 9600, 10500, 10800, 11400, 11700, 13200, 15000, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 3900, 4200, 
    4800, 6000, 7500, 8700, 9000, 9900, 10200, 10500, 11400, 12600, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7200, 9000, 10500, 15000, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    6300, 7500, 8700, 9000, 10200, 10500, 12900, 15000, 15900, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7200, 7500, 7800, 8400, 9000, 9900, 10500, 11100, 12300, 14400, 14700, 
    15000, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 8700, 9000, 9600, 10500, 13500, 13800, 14400, 15000, 15300, 15600, 
    15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4500, 
    4800, 5700, 6000, 7500, 9000, 10500, 12900, 14700, 15000, 15900, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 4800, 
    6000, 7500, 9000, 9900, 10500, 11700, 14700, 15000, 15600, 15900, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3000, 3300, 3600, 
    4200, 4500, 4800, 5100, 6000, 6300, 7500, 7800, 9000, 9300, 10500, 11400, 
    12600, 12900, 13800, 14400, 15000, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 
    4800, 6000, 7500, 9000, 10500, 12300, 13800, 15000, 15300, 15900, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 10500, 15000, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5400, 
    5700, 6000, 7500, 9000, 10500, 10800, 12000, 12600, 13200, 15000, 15900, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 600, 900, 1200, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 4800, 5400, 
    6000, 7500, 9000, 10500, 12000, 14100, 15000, 15300, 15600, 15900, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5700, 
    6000, 6600, 6900, 7500, 8100, 9000, 9900, 10500, 11700, 12600, 13800, 
    14700, 15000, 15600, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 4800, 
    6000, 6300, 7500, 9000, 9300, 10500, 10800, 12000, 12900, 13500, 13800, 
    15000, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0, 600, 900, 4200, 8400, 9000, 9600, 10200, 10500, 11400, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0, 600, 900, 1200, 1800, 2100, 2400, 2700, 3300, 3600, 4200, 4800, 6000, 
    6300, 6900, 7500, 7800, 8100, 9000, 9300, 10200, 10500, 10800, 11400, 
    12000, 12600, 13200, 13500, 14100, 14400, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 3900, 4200, 
    4800, 5400, 6000, 7500, 7800, 8100, 9000, 9600, 9900, 10500, 11400, 
    12000, 12900, 13500, 15000, 15600, 15900, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 4500, 
    4800, 6000, 6600, 7500, 9000, 9300, 9900, 10500, 11100, 11700, 12300, 
    12900, 13200, 13500, 13800, 15000, 15900, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 10500, 13500, 15000, 15900, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3000, 3600, 4200, 4800, 
    5700, 6000, 6600, 7500, 9000, 10500, 11700, 13500, 13800, 14100, 14700, 
    15000, 15300, 15900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3000, 3300, 3600, 3900, 4200, 
    4500, 4800, 5100, 6000, 7500, 9000, 10200, 10500, 11100, 11400, 11700, 
    12000, 12600, 12900, 13200, 13800, 14400, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3000, 3300, 3600, 
    3900, 4200, 4500, 4800, 5100, 5400, 5700, 6000, 6600, 7200, 7800, 8400, 
    9000, 9600, 10200, 10500, 11400, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0, 300, 600, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 6000, 
    7500, 9000, 10500, 12000, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 300, 600, 1200, 1500, 1800, 2100, 2400, 2700, 3000, 3300, 3600, 3900, 
    4200, 4500, 4800, 5100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  300, 600, 900, 1200, 1500, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5400, 
    6000, 6900, 7500, 9000, 9300, 9900, 10500, 10800, 11100, 11700, 0, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 6600, 7500, 9000, 10500, 12000, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0, 900, 1200, 1800, 2100, 2400, 2700, 3600, 4200, 4800, 5700, 6000, 7500, 
    9000, 10500, 10800, 14400, 15000, 15600, 15600, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 wdSigW =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  50, 85, 85, 90, 85, 85, 90, 90, 90, 80, 65, 40, 40, 50, 65, 75, 60, 325, 
    300, 310, 345, 10, 5, 260, 265, 270, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  180, 195, 205, 210, 215, 235, 240, 235, 235, 205, 210, 225, 235, 245, 245, 
    245, 240, 255, 250, 260, 240, 260, 310, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  325, 320, 320, 10, 330, 325, 265, 285, 280, 260, 265, 270, 250, 255, 260, 
    250, 250, 245, 240, 240, 240, 230, 255, 245, 250, 255, 240, 225, 240, 
    230, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  130, 95, 210, 235, 235, 205, 145, 140, 175, 80, 75, 40, 60, 65, 65, 60, 85, 
    105, 125, 120, 170, 205, 235, 215, 215, 245, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  60, 45, 80, 110, 150, 290, 315, 330, 345, 330, 330, 335, 310, 295, 300, 
    310, 310, 315, 325, 335, 315, 330, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  90, 165, 200, 200, 200, 215, 230, 240, 245, 245, 240, 245, 245, 245, 245, 
    250, 245, 240, 240, 225, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  80, 125, 125, 130, 110, 100, 110, 130, 155, 180, 175, 175, 175, 190, 195, 
    195, 190, 200, 200, 195, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  140, 140, 140, 150, 155, 175, 175, 180, 180, 175, 170, 165, 165, 180, 180, 
    185, 180, 180, 175, 180, 180, 190, 200, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  250, 265, 25, 85, 115, 180, 195, 200, 205, 235, 230, 235, 240, 245, 250, 
    250, 260, 265, 245, 250, 255, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  320, 315, 245, 230, 245, 230, 235, 240, 245, 245, 245, 255, 250, 250, 250, 
    255, 275, 280, 280, 255, 260, 275, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  190, 190, 195, 195, 190, 195, 210, 220, 225, 235, 245, 245, 250, 245, 260, 
    255, 250, 280, 280, 275, 255, 245, 260, 265, 280, 265, 255, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  170, 145, 150, 155, 155, 195, 190, 175, 175, 120, 90, 60, 155, 50, 125, 
    330, 340, 360, 35, 35, 35, 40, 355, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  230, 245, 245, 240, 235, 250, 250, 245, 240, 235, 235, 235, 240, 245, 245, 
    250, 245, 240, 255, 240, 225, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  340, 50, 80, 125, 170, 225, 245, 250, 250, 235, 235, 235, 240, 245, 245, 
    240, 245, 245, 240, 235, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  300, 330, 30, 45, 330, 265, 265, 260, 260, 260, 260, 260, 265, 265, 265, 
    265, 270, 270, 265, 265, 245, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  40, 0, 270, 235, 235, 260, 255, 255, 265, 280, 285, 280, 280, 280, 280, 
    285, 285, 280, 295, 285, 280, 295, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  150, 245, 320, 340, 355, 5, 10, 335, 285, 280, 280, 270, 275, 275, 275, 
    275, 275, 275, 280, 280, 275, 275, 280, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  140, 150, 225, 345, 10, 315, 305, 305, 300, 290, 295, 300, 300, 300, 305, 
    300, 305, 305, 300, 310, 325, 320, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  340, 350, 355, 15, 5, 350, 345, 350, 330, 325, 335, 340, 335, 330, 330, 
    325, 325, 330, 335, 325, 325, 330, 340, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  200, 335, 300, 240, 180, 180, 190, 195, 205, 255, 255, 260, 250, 280, 290, 
    295, 265, 245, 210, 270, 255, 310, 315, 225, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  30, 25, 5, 360, 345, 340, 15, 30, 85, 90, 85, 80, 85, 70, 75, 115, 115, 
    115, 120, 125, 130, 175, 195, 215, 210, 225, 250, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  100, 125, 140, 95, 65, 65, 65, 45, 35, 30, 50, 70, 80, 75, 50, 55, 40, 45, 
    350, 355, 295, 295, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  85, 85, 90, 95, 120, 215, 235, 235, 240, 225, 215, 220, 220, 225, 230, 240, 
    250, 235, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  350, 10, 40, 40, 360, 360, 355, 340, 335, 330, 305, 280, 280, 270, 265, 
    260, 250, 250, 255, 255, 250, 245, 260, 265, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  120, 80, 75, 60, 45, 50, 55, 60, 60, 70, 70, 70, 350, 360, 360, 355, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  330, 350, 355, 360, 355, 355, 340, 325, 315, 300, 290, 270, 260, 250, 255, 
    245, 250, 250, 250, 240, 265, 260, 235, 230, 240, 220, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  355, 10, 10, 5, 5, 5, 5, 5, 5, 10, 5, 5, 10, 40, 65, 60, 35, 25, 20, 20, 
    360, 5, 340, 10, 30, 45, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  90, 90, 90, 90, 85, 60, 55, 60, 65, 70, 55, 40, 20, 25, 55, 20, 45, 45, 25, 
    275, 275, 290, 265, 285, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0, 240, 235, 195, 195, 205, 205, 205, 165, 80, 70, 65, 60, 60, 5, 10, 25, 
    35, 60, 60, 20, 40, 65, 10, 25, 35, 330, 330, 340, 305, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  240, 265, 270, 295, 295, 290, 290, 275, 275, 300, 315, 310, 310, 310, 325, 
    30, 20, 345, 350, 360, 360, 325, 320, 310, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 305, 295, 305, 280, 265, 270, 295, 295, 300, 295, 315, 355, 330, 325, 
    335, 345, 10, 360, 335, 335, 305, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  185, 205, 230, 250, 265, 275, 265, 250, 255, 270, 310, 310, 330, 345, 340, 
    345, 20, 15, 10, 330, 315, 270, 270, 350, 320, 325, 330, 300, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  60, 90, 85, 60, 330, 305, 295, 295, 300, 295, 295, 290, 295, 315, 290, 310, 
    315, 335, 355, 345, 325, 315, 335, 300, 310, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  210, 245, 255, 250, 245, 245, 245, 255, 270, 275, 280, 285, 300, 315, 300, 
    285, 290, 300, 295, 290, 320, 310, 315, 285, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  175, 175, 180, 175, 160, 145, 195, 245, 240, 235, 240, 290, 300, 305, 290, 
    295, 300, 300, 310, 315, 335, 335, 330, 340, 325, 310, 300, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  155, 205, 225, 230, 250, 265, 265, 265, 260, 255, 255, 265, 265, 265, 295, 
    285, 300, 300, 310, 330, 315, 320, 325, 305, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  230, 240, 250, 260, 260, 250, 245, 250, 255, 245, 255, 260, 270, 275, 260, 
    265, 270, 275, 280, 290, 285, 295, 305, 290, 285, 275, 285, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 230, 260, 290, 285, 290, 290, 300, 305, 300, 315, 315, 310, 320, 325, 
    325, 315, 310, 300, 290, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  340, 70, 140, 145, 145, 235, 265, 280, 295, 355, 335, 335, 335, 325, 310, 
    310, 315, 325, 330, 330, 335, 300, 295, 300, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  350, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  190, 210, 245, 260, 265, 265, 275, 285, 280, 260, 260, 270, 280, 290, 295, 
    290, 285, 285, 265, 285, 285, 275, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  120, 185, 195, 185, 175, 145, 150, 145, 125, 65, 75, 70, 70, 60, 75, 50, 
    45, 60, 70, 35, 55, 350, 335, 325, 335, 355, 325, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  170, 175, 190, 200, 200, 195, 175, 160, 140, 130, 110, 110, 25, 235, 230, 
    265, 280, 220, 225, 275, 300, 305, 295, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  135, 155, 160, 170, 165, 160, 170, 290, 230, 290, 195, 165, 250, 275, 280, 
    290, 300, 280, 290, 290, 290, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  150, 155, 170, 185, 185, 170, 165, 145, 140, 170, 170, 195, 185, 185, 205, 
    220, 245, 235, 240, 240, 270, 280, 275, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  210, 220, 235, 235, 230, 225, 220, 205, 200, 20, 25, 45, 35, 30, 305, 290, 
    315, 290, 250, 285, 295, 315, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  190, 205, 220, 220, 220, 215, 200, 190, 185, 150, 140, 135, 145, 250, 245, 
    265, 270, 240, 225, 230, 240, 230, 275, 285, 285, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  235, 230, 220, 210, 205, 195, 190, 180, 185, 200, 240, 215, 185, 200, 205, 
    215, 230, 235, 225, 260, 265, 280, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  150, 215, 245, 260, 265, 165, 170, 185, 210, 220, 230, 235, 230, 250, 245, 
    225, 230, 250, 255, 260, 235, 255, 250, 240, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  220, 205, 200, 210, 235, 205, 195, 205, 215, 215, 225, 230, 220, 215, 225, 
    230, 230, 225, 250, 245, 250, 235, 245, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  220, 205, 215, 205, 215, 210, 215, 215, 215, 220, 225, 230, 235, 230, 220, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  190, 205, 170, 175, 185, 185, 190, 195, 195, 200, 210, 210, 210, 210, 210, 
    215, 225, 240, 220, 230, 235, 225, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  180, 225, 245, 250, 255, 260, 265, 270, 280, 290, 280, 295, 290, 320, 290, 
    240, 230, 275, 285, 300, 240, 235, 275, 280, 290, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  190, 200, 220, 225, 225, 230, 235, 245, 265, 255, 205, 220, 235, 235, 245, 
    235, 220, 220, 245, 270, 275, 280, 260, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  10, 20, 50, 75, 85, 195, 215, 225, 225, 240, 235, 225, 220, 220, 250, 265, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  130, 165, 205, 230, 235, 230, 220, 195, 185, 210, 230, 225, 225, 225, 230, 
    225, 230, 230, 265, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  210, 225, 260, 300, 300, 285, 285, 300, 300, 255, 265, 270, 250, 240, 225, 
    240, 260, 260, 255, 245, 265, 240, 260, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  340, 20, 15, 15, 310, 230, 240, 260, 260, 250, 250, 250, 255, 255, 240, 
    240, 250, 245, 245, 260, 250, 270, 270, 245, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  360, 5, 20, 40, 35, 35, 100, 175, 210, 225, 230, 240, 240, 240, 240, 240, 
    240, 230, 240, 265, 255, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  130, 15, 55, 70, 180, 200, 200, 200, 205, 210, 210, 220, 215, 235, 230, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  240, 245, 265, 285, 285, 285, 280, 275, 280, 285, 285, 275, 275, 280, 280, 
    280, 260, 255, 250, 275, 275, 270, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  360, 15, 15, 5, 325, 320, 330, 340, 335, 310, 295, 290, 285, 280, 275, 270, 
    255, 255, 255, 255, 250, 250, 270, 260, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  100, 80, 310, 270, 225, 210, 215, 210, 230, 240, 225, 215, 220, 215, 210, 
    215, 215, 210, 210, 230, 235, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  330, 345, 360, 360, 360, 355, 350, 350, 320, 305, 290, 285, 275, 265, 260, 
    265, 275, 270, 265, 255, 270, 270, 270, 265, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  90, 110, 115, 210, 335, 350, 345, 280, 265, 285, 265, 270, 270, 250, 250, 
    250, 245, 245, 250, 260, 260, 260, 35, 360, 290, 290, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  10, 25, 50, 130, 90, 50, 45, 5, 355, 40, 90, 75, 40, 95, 20, 30, 30, 55, 
    250, 280, 270, 275, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  80, 90, 100, 95, 80, 80, 100, 90, 60, 5, 340, 340, 330, 305, 5, 305, 300, 
    285, 290, 280, 330, 360, 5, 10, 35, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  360, 75, 80, 80, 85, 85, 100, 95, 90, 85, 85, 75, 90, 75, 65, 80, 70, 85, 
    100, 95, 90, 95, 90, 70, 75, 80, 90, 75, 70, 85, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 175, 130, 55, 30, 35, 30, 25, 335, 330, 345, 355, 355, 345, 335, 330, 
    335, 340, 350, 350, 285, 295, 305, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  160, 185, 195, 195, 185, 205, 215, 215, 225, 225, 230, 235, 245, 260, 270, 
    275, 285, 295, 300, 305, 290, 305, 300, 285, 295, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  210, 280, 320, 325, 335, 330, 335, 325, 315, 320, 325, 320, 320, 320, 320, 
    320, 315, 315, 310, 285, 290, 295, 270, 280, 275, 265, 240, 255, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  150, 165, 180, 190, 200, 250, 250, 245, 235, 260, 275, 280, 285, 275, 275, 
    280, 280, 285, 285, 290, 285, 290, 290, 275, 270, 295, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  295, 305, 280, 260, 245, 240, 240, 235, 230, 215, 215, 220, 225, 230, 225, 
    230, 230, 235, 235, 245, 255, 245, 250, 275, 265, 255, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  90, 110, 125, 130, 130, 250, 250, 255, 270, 290, 285, 280, 275, 285, 310, 
    305, 320, 320, 340, 350, 355, 325, 305, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  60, 85, 95, 90, 85, 70, 65, 70, 85, 60, 55, 45, 330, 310, 330, 285, 255, 
    265, 280, 280, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  210, 180, 195, 165, 25, 35, 40, 50, 60, 45, 20, 360, 350, 345, 360, 15, 30, 
    45, 30, 15, 45, 50, 360, 355, 325, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  210, 225, 245, 250, 230, 290, 355, 355, 40, 120, 100, 35, 5, 320, 320, 335, 
    315, 280, 315, 315, 325, 350, 320, 330, 330, 330, 20, 40, 40, 30, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 125, 125, 360, 285, 150, 30, 50, 75, 355, 360, 35, 45, 45, 355, 340, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  270, 275, 290, 300, 300, 280, 280, 270, 280, 15, 30, 30, 30, 340, 45, 35, 
    35, 30, 25, 60, 40, 355, 355, 345, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  190, 180, 185, 175, 175, 170, 170, 175, 170, 140, 140, 115, 90, 80, 60, 30, 
    45, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  180, 205, 215, 205, 200, 190, 185, 185, 155, 120, 110, 105, 100, 100, 105, 
    105, 35, 35, 30, 20, 55, 290, 265, 285, 310, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 290, 310, 310, 295, 290, 285, 285, 285, 280, 295, 300, 285, 290, 335, 
    325, 330, 335, 315, 310, 305, 345, 345, 15, 360, 335, 335, 310, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  360, 55, 100, 105, 105, 100, 50, 325, 310, 315, 305, 295, 310, 315, 315, 
    305, 300, 300, 310, 310, 320, 340, 310, 310, 305, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  160, 235, 230, 240, 245, 245, 255, 250, 250, 245, 250, 275, 290, 300, 310, 
    305, 315, 320, 300, 300, 300, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  130, 95, 95, 95, 95, 90, 100, 110, 115, 190, 260, 275, 265, 250, 255, 255, 
    275, 270, 275, 260, 255, 265, 260, 270, 280, 285, 330, 305, 325, 300, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  140, 150, 160, 160, 160, 150, 145, 150, 125, 110, 40, 340, 25, 15, 330, 
    305, 300, 310, 315, 310, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  140, 150, 155, 160, 160, 160, 155, 170, 170, 110, 60, 10, 30, 10, 15, 15, 
    315, 310, 300, 305, 310, 310, 310, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  110, 125, 190, 220, 220, 235, 235, 230, 220, 210, 200, 205, 225, 230, 230, 
    235, 235, 245, 250, 235, 245, 235, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  260, 235, 195, 215, 265, 255, 255, 255, 250, 240, 235, 240, 230, 230, 225, 
    225, 230, 235, 240, 240, 235, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  300, 230, 155, 100, 110, 180, 195, 195, 200, 215, 225, 225, 215, 215, 220, 
    235, 215, 230, 255, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  140, 175, 180, 185, 190, 200, 200, 200, 195, 205, 210, 215, 215, 215, 225, 
    220, 240, 230, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 115, 200, 235, 40, 75, 95, 85, 35, 30, 40, 50, 50, 35, 40, 40, 30, 30, 
    265, 245, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  200, 220, 235, 235, 245, 250, 250, 250, 250, 250, 260, 265, 270, 280, 280, 
    280, 290, 265, 265, 270, 265, 295, 270, 280, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  290, 290, 305, 315, 295, 270, 275, 275, 265, 265, 270, 265, 260, 270, 265, 
    260, 255, 255, 255, 255, 270, 260, 250, 250, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  340, 15, 25, 35, 335, 275, 245, 255, 265, 245, 240, 250, 240, 240, 260, 
    265, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  210, 200, 125, 140, 140, 125, 115, 135, 180, 230, 230, 230, 225, 215, 230, 
    230, 230, 245, 230, 250, 255, 250, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 335, 320, 360, 20, 30, 10, 360, 5, 10, 355, 360, 25, 20, 10, 25, 20, 20, 
    20, 20, 25, 20, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  220, 225, 240, 265, 275, 270, 265, 270, 285, 295, 280, 275, 275, 275, 270, 
    260, 270, 270, 280, 265, 260, 280, 20, 5, 360, 355, 340, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 125, 145, 140, 135, 130, 140, 135, 125, 85, 105, 100, 95, 330, 300, 280, 
    215, 185, 230, 220, 260, 290, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  160, 0, 315, 280, 225, 170, 130, 120, 115, 120, 120, 120, 90, 95, 155, 50, 
    40, 30, 5, 360, 360, 340, 10, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  60, 65, 70, 75, 85, 95, 105, 115, 135, 120, 110, 130, 150, 60, 300, 240, 
    280, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  40, 25, 45, 50, 60, 65, 60, 60, 55, 25, 25, 25, 20, 20, 25, 5, 10, 25, 25, 
    5, 15, 30, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  90, 165, 180, 195, 250, 280, 295, 315, 320, 320, 315, 305, 310, 300, 305, 
    305, 305, 310, 320, 315, 315, 310, 305, 295, 290, 280, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  230, 285, 285, 280, 270, 310, 315, 310, 310, 310, 315, 320, 325, 325, 325, 
    325, 325, 315, 295, 280, 290, 265, 275, 275, 260, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  340, 350, 340, 355, 350, 300, 300, 295, 295, 280, 285, 285, 290, 285, 275, 
    275, 270, 270, 270, 260, 280, 275, 270, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  330, 335, 350, 350, 335, 320, 315, 310, 310, 305, 300, 300, 300, 290, 285, 
    285, 275, 280, 285, 275, 275, 285, 270, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  120, 145, 145, 145, 140, 135, 140, 155, 160, 165, 170, 200, 200, 250, 255, 
    260, 270, 260, 255, 270, 270, 265, 255, 245, 240, 205, 195, 190, 170, 
    175, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  280, 330, 25, 65, 70, 60, 55, 55, 50, 60, 75, 75, 70, 70, 75, 70, 70, 80, 
    80, 55, 75, 75, 55, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  60, 110, 80, 350, 330, 335, 335, 330, 325, 325, 330, 330, 325, 315, 310, 
    310, 320, 325, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 310, 330, 330, 330, 330, 325, 330, 325, 320, 315, 305, 315, 320, 320, 
    315, 310, 310, 310, 310, 325, 310, 330, 320, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  240, 300, 350, 345, 340, 350, 350, 330, 300, 315, 300, 305, 300, 305, 310, 
    315, 310, 305, 325, 320, 305, 330, 330, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  290, 310, 310, 310, 310, 315, 325, 325, 320, 325, 330, 325, 320, 320, 315, 
    315, 315, 305, 315, 325, 320, 315, 330, 320, 325, 335, 350, 340, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 230, 245, 240, 230, 230, 225, 230, 225, 240, 250, 245, 240, 250, 255, 
    255, 255, 255, 255, 255, 260, 275, 270, 265, 270, 280, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  110, 295, 355, 255, 120, 210, 210, 240, 250, 270, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  90, 185, 205, 170, 260, 325, 15, 335, 345, 360, 10, 315, 310, 305, 330, 
    305, 325, 315, 325, 335, 315, 320, 335, 325, 330, 305, 325, 315, 335, 
    290, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  350, 10, 15, 10, 5, 360, 350, 335, 330, 320, 330, 330, 320, 305, 280, 285, 
    275, 275, 270, 255, 250, 245, 255, 260, 260, 280, 265, 295, 290, 265, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  230, 315, 30, 45, 55, 55, 55, 55, 50, 50, 70, 55, 50, 55, 55, 40, 55, 45, 
    45, 55, 30, 40, 15, 45, 20, 60, 25, 10, 75, 50, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  310, 335, 335, 335, 335, 335, 335, 335, 330, 340, 355, 355, 360, 360, 360, 
    15, 30, 70, 85, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  245, 300, 290, 335, 330, 310, 295, 305, 320, 330, 340, 350, 5, 350, 350, 
    345, 350, 355, 355, 355, 355, 335, 325, 335, 350, 10, 345, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  30, 65, 75, 60, 40, 360, 355, 340, 320, 325, 310, 285, 300, 295, 295, 285, 
    305, 280, 275, 275, 285, 290, 280, 295, 270, 280, 300, 275, 300, 270, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 105, 85, 80, 80, 80, 80, 90, 90, 110, 115, 125, 125, 95, 80, 75, 55, 55, 
    70, 90, 105, 255, 265, 260, 250, 250, 265, 290, 315, 285, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  260, 280, 290, 275, 260, 205, 200, 205, 205, 225, 215, 220, 220, 225, 220, 
    230, 235, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  10, 45, 75, 105, 95, 115, 110, 110, 130, 135, 160, 205, 240, 275, 300, 325, 
    105, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  115, 115, 110, 110, 100, 105, 110, 70, 90, 85, 110, 95, 110, 95, 90, 95, 
    110, 110, 105, 155, 145, 145, 165, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  310, 250, 255, 250, 235, 240, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  210, 235, 260, 295, 300, 280, 275, 280, 250, 245, 230, 230, 225, 225, 225, 
    225, 235, 245, 240, 240, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 wsSigW =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  3, 8.7, 8.2, 8.7, 8.7, 8.2, 8.7, 9.2, 10.2, 7.7, 5.6, 5.6, 5.1, 3.6, 3.6, 
    3.6, 2, 3, 2.5, 2.5, 1.5, 2.5, 0.5, 2.5, 6.6, 26.7, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 5.6, 6.1, 5.6, 5.6, 6.1, 6.6, 8.2, 7.7, 7.2, 8.2, 8.7, 8.2, 8.2, 9.7, 
    13.3, 15.4, 12.3, 9.2, 7.2, 6.1, 4.6, 3, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  4.1, 11.8, 11.3, 5.6, 3, 0.5, 5.1, 7.2, 8.7, 10.2, 8.7, 7.7, 7.2, 13.3, 
    17.5, 20, 23.6, 22.6, 24.1, 32.4, 27.2, 26.2, 26.2, 19.5, 25.2, 20.5, 19, 
    22.1, 22.1, 22.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  2, 0.5, 0.5, 1.5, 2.5, 2, 1.5, 2, 1.5, 3.6, 4.6, 7.2, 8.7, 8.2, 6.6, 6.1, 
    4.6, 6.1, 8.7, 7.2, 5.6, 6.6, 10.2, 14.4, 13.8, 12.8, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 2.5, 4.6, 3.6, 2.5, 2.5, 5.1, 7.7, 7.7, 7.2, 8.7, 7.7, 8.7, 12.3, 
    12.8, 18, 21.6, 23.1, 22.6, 9.7, 11.8, 9.7, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 5.1, 6.1, 7.2, 9.2, 8.7, 9.7, 10.2, 11.3, 13.8, 17.5, 20.5, 24.1, 41.6, 
    53.5, 57.1, 40.1, 31.9, 5.6, 9.2, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6.6, 12.3, 11.8, 11.3, 11.3, 12.3, 11.3, 11.3, 11.8, 13.8, 19, 21.6, 21.6, 
    25.7, 26.2, 29.3, 40.6, 16.4, 10.8, 8.7, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  10.2, 13.3, 15.9, 15.4, 11.3, 3.6, 3, 4.1, 7.7, 11.8, 11.8, 11.3, 11.3, 
    13.8, 14.4, 16.4, 16.9, 16.9, 21.6, 28.8, 13.8, 12.8, 6.6, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 1.5, 1, 2.5, 3, 4.6, 5.6, 5.6, 5.6, 7.7, 9.7, 14.4, 13.8, 14.9, 18, 
    22.6, 26.2, 25.2, 12.3, 12.3, 6.6, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.6, 1.5, 1.5, 3, 4.1, 7.2, 7.7, 7.2, 6.6, 8.2, 9.2, 12.8, 13.8, 15.4, 
    15.9, 16.4, 17.5, 16.9, 23.1, 13.3, 12.3, 5.6, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.1, 3.6, 4.6, 7.2, 9.2, 9.2, 9.2, 11.3, 11.8, 11.3, 12.3, 10.8, 9.2, 10.8, 
    11.3, 9.7, 9.7, 11.3, 12.8, 10.2, 13.3, 13.3, 9.7, 15.9, 14.4, 10.2, 5.1, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2.5, 2.5, 1, 1.5, 2, 2.5, 3.6, 3.6, 2, 2.5, 1.5, 3.6, 5.1, 6.6, 
    8.7, 22.6, 29.3, 24.1, 20.5, 5.6, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  2.5, 9.7, 9.7, 9.2, 8.7, 12.3, 12.8, 12.8, 12.3, 11.3, 10.2, 13.3, 21.1, 
    28.8, 33.4, 32.9, 29.8, 22.1, 16.9, 7.2, 8.2, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 6.6, 4.6, 2.5, 3, 4.1, 4.1, 6.6, 7.2, 9.7, 11.8, 13.8, 23.1, 26.7, 33.4, 
    38.6, 42.2, 23.1, 13.8, 9.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1.5, 0.5, 1, 1, 5.1, 5.6, 5.6, 6.1, 8.2, 13.3, 18.5, 19.5, 25.7, 38.6, 
    41.6, 46.3, 48.3, 23.6, 10.8, 7.7, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5, 0, 0.5, 2, 3, 3, 3.6, 4.6, 8.7, 12.8, 13.8, 12.8, 16.4, 22.1, 25.7, 
    31.4, 26.7, 22.1, 14.4, 9.7, 10.2, 9.7, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3.6, 3.6, 3, 5.6, 5.6, 6.1, 5.1, 7.2, 10.2, 10.2, 13.8, 16.9, 23.1, 
    24.7, 27.2, 25.7, 31.9, 43.2, 33.4, 19.5, 14.9, 10.8, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 1, 2.5, 1, 4.1, 6.1, 7.2, 9.2, 10.8, 12.3, 15.9, 19, 25.7, 28.3, 
    33.9, 38.6, 41.1, 16.9, 14.9, 9.7, 9.7, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 7.2, 5.1, 3, 2.5, 4.1, 4.1, 5.1, 6.1, 8.7, 11.8, 13.3, 14.4, 19, 23.1, 
    24.1, 26.7, 33.4, 32.9, 38.6, 14.9, 13.8, 10.8, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.5, 2.5, 1.5, 1.5, 5.6, 5.1, 5.6, 5.6, 5.1, 7.2, 7.7, 7.2, 6.6, 6.6, 6.6, 
    7.2, 8.7, 8.7, 9.2, 6.6, 9.2, 6.6, 7.2, 4.6, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 5.1, 5.6, 4.1, 3, 2, 2, 1.5, 1.5, 5.6, 6.1, 8.7, 10.2, 10.8, 10.8, 
    7.2, 5.6, 8.2, 11.8, 11.3, 9.7, 8.2, 9.7, 9.2, 21.1, 17.5, 13.3, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4.6, 3.6, 2, 4.1, 5.6, 4.1, 4.1, 5.1, 5.6, 6.1, 4.1, 2.5, 2, 3.6, 7.7, 
    10.2, 7.7, 7.7, 8.2, 6.6, 8.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.6, 6.1, 7.2, 5.6, 3, 9.2, 10.8, 11.8, 16.9, 21.6, 28.3, 35, 42.2, 46.3, 
    21.1, 20, 15.9, 9.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4.6, 9.2, 9.2, 9.7, 8.7, 7.7, 8.7, 10.2, 9.2, 9.2, 12.3, 14.4, 24.7, 
    28.8, 36, 37, 36.5, 43.7, 47.8, 46.3, 31.4, 18.5, 13.3, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.5, 5.1, 5.6, 6.6, 6.6, 6.6, 6.6, 6.6, 6.6, 8.2, 6.1, 3.6, 2, 5.6, 6.6, 
    5.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.6, 7.7, 12.8, 13.8, 11.8, 13.8, 13.3, 11.8, 12.8, 12.8, 14.4, 16.4, 24.7, 
    26.7, 29.3, 36.5, 48.3, 40.6, 24.1, 23.1, 19.5, 12.3, 9.7, 10.2, 10.2, 
    10.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  12.3, 12.3, 11.8, 11.3, 11.3, 12.3, 12.8, 13.3, 12.8, 12.8, 12.3, 12.3, 
    11.8, 9.2, 9.2, 9.2, 10.2, 9.2, 7.2, 7.2, 5.6, 5.6, 5.6, 5.6, 6.6, 6.1, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1, 7.7, 7.7, 7.7, 7.7, 7.2, 7.7, 7.7, 7.7, 7.2, 5.1, 4.6, 5.6, 5.1, 3, 3.6, 
    4.6, 6.1, 4.6, 7.2, 15.9, 14.4, 10.8, 9.7, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 10.8, 8.7, 9.2, 9.2, 5.6, 5.6, 4.6, 3, 6.1, 6.6, 8.7, 10.2, 6.6, 4.6, 
    7.2, 8.2, 6.1, 5.6, 7.7, 7.2, 7.2, 7.2, 10.8, 11.8, 8.7, 10.2, 10.2, 7.2, 
    5.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 12.3, 10.8, 7.7, 6.6, 3.6, 4.1, 4.1, 4.6, 5.6, 6.1, 6.1, 5.6, 7.2, 4.6, 
    4.6, 5.6, 7.7, 7.7, 12.3, 16.9, 8.7, 8.7, 8.2, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 5.6, 6.1, 5.1, 4.6, 5.6, 6.1, 7.2, 6.6, 6.1, 5.6, 5.1, 6.6, 6.1, 10.8, 
    12.3, 13.3, 17.5, 21.1, 11.8, 9.7, 6.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 6.6, 13.3, 11.8, 11.8, 12.3, 9.7, 9.2, 9.2, 8.7, 7.2, 8.7, 12.3, 10.2, 
    7.2, 7.2, 8.7, 9.2, 7.2, 7.2, 9.2, 7.2, 6.1, 6.1, 5.6, 9.2, 7.2, 6.6, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7.2, 6.1, 6.6, 3.6, 3.6, 6.6, 7.2, 6.6, 5.6, 6.6, 7.7, 7.2, 6.6, 6.6, 10.8, 
    16.9, 16.9, 20, 30.8, 23.1, 8.7, 11.8, 10.8, 10.2, 13.3, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.6, 14.4, 14.9, 14.4, 13.8, 13.8, 12.8, 11.8, 11.8, 10.2, 10.8, 9.2, 6.6, 
    9.7, 11.8, 9.7, 10.2, 14.4, 13.8, 14.4, 23.6, 10.8, 7.2, 7.2, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.5, 4.1, 6.1, 6.6, 6.1, 4.1, 3, 2.5, 3, 4.6, 5.1, 4.1, 7.7, 10.8, 14.9, 
    15.4, 15.4, 19.5, 20.5, 25.2, 40.1, 32.4, 37.5, 23.1, 17.5, 14.4, 13.8, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 8.7, 8.7, 9.2, 8.7, 10.8, 11.8, 13.3, 14.4, 14.9, 10.2, 9.7, 10.8, 10.8, 
    11.8, 14.9, 12.3, 12.8, 22.1, 29.3, 20, 14.4, 12.3, 8.7, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.1, 16.4, 16.4, 18.5, 20, 18.5, 17.5, 15.4, 16.4, 14.4, 12.3, 13.8, 16.4, 
    16.9, 18.5, 22.1, 25.2, 20.5, 16.9, 20.5, 21.6, 40.6, 29.8, 13.3, 10.2, 
    11.8, 10.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 2.5, 2, 5.6, 7.2, 8.2, 7.7, 12.3, 10.8, 12.8, 14.9, 15.4, 24.7, 30.3, 
    36.5, 38.6, 39.1, 24.7, 16.4, 13.8, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.5, 3.6, 4.6, 4.1, 3, 1.5, 2.5, 3, 3.6, 2.5, 4.6, 8.2, 12.3, 17.5, 17.5, 
    20, 19.5, 23.6, 29.3, 30.3, 23.1, 13.8, 14.4, 19, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  3.6, 9.7, 19.5, 18.5, 15.4, 9.7, 10.8, 12.3, 14.4, 15.4, 15.4, 13.3, 14.9, 
    13.3, 13.3, 15.9, 14.4, 13.3, 20, 15.4, 11.8, 10.8, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5, 4.1, 4.1, 4.6, 5.6, 4.6, 5.1, 4.1, 2, 3.6, 5.6, 8.2, 7.2, 4.1, 4.1, 
    6.1, 7.7, 14.9, 11.8, 13.3, 7.7, 6.6, 8.7, 9.2, 8.2, 6.1, 7.7, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.1, 6.6, 11.8, 13.3, 13.3, 9.2, 9.2, 10.8, 13.8, 11.8, 10.8, 7.7, 1.5, 
    4.1, 4.1, 5.6, 6.1, 6.6, 7.7, 13.8, 14.9, 14.4, 14.9, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.6, 13.8, 13.8, 12.8, 11.8, 10.2, 5.6, 1, 2.5, 3.6, 2, 8.2, 9.2, 12.3, 
    14.9, 24.1, 21.1, 21.6, 26.2, 24.1, 13.3, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.6, 6.1, 14.9, 12.8, 7.7, 5.6, 5.1, 4.6, 3.6, 5.1, 5.6, 5.6, 7.2, 9.7, 
    12.8, 10.2, 6.1, 8.2, 12.8, 12.8, 22.1, 18.5, 15.4, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 7.7, 16.4, 15.9, 13.8, 10.2, 8.2, 6.1, 5.1, 2.5, 5.1, 3.6, 5.1, 4.1, 
    2, 6.6, 7.7, 6.1, 7.2, 12.8, 11.8, 4.6, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.1, 21.1, 19.5, 15.9, 9.7, 9.2, 9.2, 9.7, 9.2, 9.2, 9.7, 7.2, 5.1, 4.1, 
    8.2, 8.7, 7.2, 7.2, 8.2, 8.2, 10.2, 10.8, 15.9, 15.9, 12.3, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.6, 8.7, 15.9, 15.4, 14.4, 14.4, 14.4, 13.3, 10.2, 8.2, 5.6, 2.5, 7.2, 
    11.3, 10.8, 13.8, 13.8, 15.4, 14.9, 23.1, 19.5, 18, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 6.6, 5.6, 5.1, 3.6, 1, 5.1, 6.1, 9.7, 12.8, 13.3, 20.5, 16.4, 17.5, 
    18, 17.5, 16.9, 16.9, 32.4, 25.2, 25.2, 26.7, 23.1, 16.4, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 6.6, 7.2, 4.1, 2, 8.2, 9.7, 11.3, 15.4, 18.5, 20.5, 19, 16.4, 16.4, 
    17.5, 17.5, 22.6, 28.3, 22.6, 27.7, 20, 15.4, 21.6, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 8.2, 9.7, 16.9, 16.4, 19.5, 21.1, 19.5, 23.1, 20, 27.7, 40.1, 28.8, 
    22.6, 16.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.5, 3.6, 4.6, 7.7, 9.7, 11.3, 14.4, 11.8, 9.2, 9.7, 13.8, 20, 31.4, 37.5, 
    43.2, 43.2, 40.1, 14.4, 18.5, 24.7, 24.1, 12.3, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 19, 21.6, 23.6, 19.5, 16.9, 15.9, 13.3, 10.8, 7.2, 6.6, 5.1, 7.2, 6.1, 
    5.6, 4.1, 3.6, 5.6, 8.7, 7.7, 8.2, 7.7, 14.4, 14.4, 5.6, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.6, 11.3, 22.1, 22.1, 21.6, 20.5, 20.5, 20, 16.9, 10.8, 7.7, 9.2, 14.9, 
    15.4, 16.9, 19, 19, 20.5, 24.1, 15.9, 14.4, 10.8, 9.7, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2.5, 2.5, 4.1, 5.6, 3, 12.3, 16.4, 24.1, 18, 18, 18, 25.2, 34.4, 22.1, 
    15.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.1, 5.1, 5.6, 7.7, 8.2, 7.2, 7.2, 8.2, 10.8, 21.1, 25.7, 30.3, 29.8, 30.3, 
    25.7, 34.4, 25.2, 25.2, 19.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 4.6, 3.6, 5.1, 3.6, 3, 4.1, 3, 3.6, 6.1, 5.6, 5.1, 5.6, 3.6, 5.6, 6.1, 
    17.5, 18, 15.9, 14.9, 12.8, 11.8, 12.8, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 6.6, 5.6, 2.5, 2, 3, 6.6, 13.3, 14.9, 17.5, 19, 19, 20, 20.5, 21.6, 
    22.1, 24.1, 31.9, 31.4, 27.2, 23.1, 13.8, 10.8, 9.2, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 6.1, 16.4, 12.3, 7.2, 5.6, 3.6, 7.2, 12.8, 16.4, 16.9, 20.5, 23.1, 
    26.7, 28.3, 25.7, 27.2, 28.8, 20.5, 22.6, 15.4, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 1, 5.6, 9.2, 15.9, 23.6, 32.4, 34.4, 36.5, 18, 22.6, 16.4, 10.8, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 5.1, 11.3, 13.8, 16.9, 16.4, 14.4, 13.8, 13.3, 13.8, 18, 23.6, 28.3, 
    34.4, 31.9, 31.9, 33.4, 30.3, 31.4, 34.4, 14.9, 13.8, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.7, 19, 17.5, 14.9, 10.8, 10.8, 10.2, 12.3, 12.3, 12.8, 18, 19, 21.6, 
    24.7, 25.2, 30.8, 37.5, 33.9, 39.1, 46.8, 49.9, 30.8, 23.1, 14.9, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2, 2, 2.5, 3.6, 4.1, 4.1, 3, 6.6, 7.7, 8.7, 8.2, 10.8, 14.4, 15.9, 14.9, 
    21.1, 26.7, 22.6, 16.4, 10.8, 10.8, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.6, 12.8, 13.3, 12.8, 11.8, 12.8, 12.3, 13.8, 13.3, 16.9, 19.5, 21.6, 
    26.2, 30.3, 29.8, 43.7, 55.5, 47.3, 47.3, 45.3, 43.2, 30.3, 21.6, 13.8, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.5, 4.1, 4.1, 1, 2, 3.6, 2.5, 6.6, 9.7, 7.2, 7.7, 8.2, 8.7, 11.8, 33.9, 
    39.1, 45.3, 49.9, 21.1, 24.1, 19.5, 13.3, 7.2, 6.6, 4.1, 3.6, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 3, 3, 2.5, 4.1, 4.1, 1.5, 4.1, 1.5, 1.5, 6.6, 2, 2.5, 7.7, 6.1, 6.1, 
    7.7, 5.6, 5.6, 6.6, 7.7, 6.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.6, 7.2, 7.2, 6.1, 4.6, 3, 3, 3, 2.5, 1.5, 3, 4.6, 6.1, 5.1, 5.6, 7.7, 
    5.6, 6.1, 6.6, 7.2, 7.7, 13.8, 17.5, 16.9, 9.7, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 9.2, 8.2, 7.2, 6.6, 6.6, 7.2, 6.6, 6.1, 6.6, 9.2, 11.3, 11.3, 13.8, 
    14.4, 16.9, 18.5, 13.3, 9.7, 9.2, 9.2, 7.7, 8.7, 9.7, 9.2, 8.2, 6.1, 7.7, 
    7.7, 6.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 4.1, 4.1, 3, 4.1, 4.6, 7.2, 6.6, 6.1, 7.7, 10.2, 12.8, 13.3, 13.8, 13.8, 
    16.9, 22.6, 26.2, 30.3, 28.8, 17.5, 18.5, 11.8, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 8.2, 10.8, 12.3, 13.3, 12.8, 14.4, 14.9, 14.4, 12.3, 13.3, 15.9, 16.4, 
    19, 20, 22.6, 20.5, 26.2, 44.2, 51.4, 25.2, 19.5, 16.4, 15.4, 16.4, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2.5, 5.6, 8.7, 9.2, 13.8, 13.8, 13.3, 12.3, 13.3, 14.4, 14.9, 18.5, 
    23.6, 28.8, 26.7, 30.3, 32.4, 27.2, 26.2, 29.3, 25.2, 20, 16.9, 13.3, 
    10.8, 12.3, 11.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  5.1, 10.2, 12.8, 12.8, 13.3, 12.3, 10.8, 11.3, 14.4, 18, 19.5, 21.6, 21.6, 
    26.2, 27.7, 28.3, 27.7, 26.7, 29.3, 37, 33.4, 16.4, 11.3, 8.2, 7.2, 4.6, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  7.7, 8.2, 6.6, 8.7, 12.8, 18, 18.5, 20.5, 21.6, 23.6, 26.2, 29.8, 31.4, 
    32.4, 31.9, 36.5, 35.5, 37.5, 31.4, 29.3, 25.7, 19, 11.3, 9.2, 7.7, 5.1, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.5, 4.6, 4.1, 3, 1.5, 4.1, 6.1, 8.2, 8.2, 8.2, 5.6, 6.1, 8.2, 8.2, 12.3, 
    13.3, 16.4, 18, 21.1, 25.7, 29.3, 11.8, 7.7, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 8.7, 9.7, 10.2, 9.7, 8.7, 8.7, 8.2, 7.2, 3.6, 4.1, 3.6, 3, 5.1, 3.6, 
    8.7, 28.8, 13.8, 12.8, 10.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.5, 6.6, 4.6, 1, 2, 4.1, 3.6, 3, 3, 4.6, 3.6, 1, 1.5, 4.6, 5.6, 4.6, 6.6, 
    5.6, 5.6, 8.7, 12.3, 10.2, 9.2, 6.6, 5.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 8.7, 7.2, 4.1, 2.5, 1, 1, 1, 1, 1, 1, 1.5, 2.5, 2.5, 2.5, 3, 3, 3.6, 
    5.1, 5.1, 4.1, 4.6, 5.1, 3.6, 4.1, 4.1, 5.1, 8.7, 8.7, 17.5, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 3, 1.5, 1, 1, 2, 2, 3.6, 2, 3.6, 5.6, 7.7, 7.7, 8.2, 6.6, 4.6, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  1, 2, 5.6, 4.6, 3.6, 2, 1.5, 1, 1.5, 4.1, 5.6, 6.1, 5.6, 2, 6.1, 5.6, 5.6, 
    9.2, 13.3, 10.8, 6.6, 6.6, 8.2, 6.1, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 7.7, 7.7, 7.7, 8.7, 8.7, 7.7, 7.7, 7.2, 7.7, 5.6, 7.7, 8.2, 6.1, 5.1, 
    5.6, 8.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 9.2, 10.8, 10.8, 9.7, 6.6, 7.2, 7.2, 7.2, 11.3, 10.2, 10.2, 10.8, 9.2, 
    6.1, 2.5, 6.6, 7.7, 6.1, 3, 0.5, 5.6, 5.6, 8.2, 14.4, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 6.6, 7.7, 8.2, 8.2, 7.2, 6.1, 7.2, 9.2, 8.7, 7.2, 6.1, 6.1, 5.6, 5.6, 
    9.2, 7.7, 7.2, 6.1, 7.7, 10.2, 12.3, 13.8, 15.4, 21.6, 11.8, 10.2, 7.7, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5, 4.1, 6.1, 7.7, 10.2, 5.6, 1, 1.5, 2.5, 3, 5.6, 6.1, 7.7, 8.7, 9.7, 
    13.8, 16.4, 19, 18.5, 22.1, 27.2, 23.6, 12.3, 12.8, 15.9, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 10.8, 9.7, 10.8, 11.8, 11.3, 11.3, 11.8, 12.3, 10.2, 13.3, 14.4, 18, 
    18.5, 24.1, 29.8, 42.2, 20.5, 21.1, 14.9, 11.3, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 9.7, 9.7, 10.2, 11.3, 8.2, 6.1, 4.1, 3.6, 2.5, 3, 7.7, 9.7, 11.8, 11.8, 
    16.4, 20.5, 24.1, 26.7, 27.7, 29.8, 33.4, 26.7, 36, 30.8, 14.9, 7.2, 7.2, 
    12.3, 7.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.6, 10.8, 11.3, 10.8, 10.8, 8.2, 7.2, 3, 2.5, 4.1, 3.6, 4.1, 5.6, 7.2, 
    8.7, 10.8, 15.4, 27.7, 24.7, 19.5, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 10.8, 11.3, 11.8, 11.8, 8.7, 5.6, 4.1, 3.6, 4.6, 4.1, 5.1, 4.6, 6.1, 
    7.2, 5.6, 4.1, 7.2, 11.8, 9.2, 25.2, 22.1, 17.5, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 1.5, 1.5, 6.1, 7.7, 9.7, 10.2, 16.4, 18, 20, 24.1, 21.1, 18.5, 19, 19, 
    29.3, 35, 44.2, 22.1, 25.7, 29.3, 19.5, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 1.5, 3.6, 8.7, 10.8, 11.8, 13.3, 15.9, 16.9, 17.5, 25.2, 33.4, 
    34.4, 35.5, 40.6, 47.8, 36.5, 25.7, 14.9, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.5, 1.5, 1, 2, 2.5, 5.6, 6.1, 6.1, 9.7, 9.2, 9.2, 10.8, 17.5, 18, 21.1, 
    18.5, 14.4, 15.9, 10.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 6.6, 8.2, 10.2, 10.2, 8.7, 11.3, 14.4, 17.5, 21.6, 29.8, 38, 40.6, 43.7, 
    34.4, 23.6, 22.6, 16.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 1.5, 1.5, 1, 2, 2.5, 2.5, 2, 4.1, 3.6, 5.6, 8.2, 9.7, 15.4, 14.9, 15.9, 
    8.7, 5.6, 4.6, 6.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.1, 26.2, 25.2, 23.6, 21.6, 21.6, 22.1, 21.6, 21.1, 18.5, 15.9, 16.9, 
    21.1, 24.1, 32.4, 30.3, 29.8, 19.5, 30.3, 26.2, 42.2, 36.5, 14.9, 14.4, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2, 2.5, 9.2, 9.7, 10.8, 14.4, 16.4, 18.5, 20, 22.6, 32.9, 34.4, 38.6, 36.5, 
    37.5, 36.5, 38, 47.3, 53.5, 49.9, 15.9, 12.3, 12.8, 17.5, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.5, 8.7, 8.2, 6.1, 2.5, 4.1, 9.2, 12.8, 14.9, 25.2, 28.3, 34.4, 36, 40.1, 
    22.1, 15.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 4.1, 4.6, 4.1, 5.6, 6.6, 7.2, 7.2, 4.1, 6.1, 7.7, 9.7, 7.7, 8.2, 21.1, 
    31.9, 31.4, 21.1, 20, 16.9, 15.9, 12.8, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 2, 3, 5.1, 7.7, 6.6, 5.6, 5.6, 6.6, 6.1, 7.7, 6.6, 5.6, 6.1, 7.2, 7.2, 
    10.2, 18.5, 23.6, 25.7, 31.9, 39.1, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6.1, 8.7, 15.9, 15.9, 15.4, 9.7, 10.2, 11.3, 12.3, 13.3, 12.8, 12.8, 14.4, 
    21.1, 21.6, 27.2, 25.2, 22.1, 21.1, 18.5, 14.4, 14.4, 9.7, 7.7, 13.3, 
    6.6, 6.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 0.5, 1, 2.5, 1.5, 2, 2, 2.5, 2.5, 3, 1.5, 3, 2, 6.6, 4.1, 5.6, 8.2, 5.6, 
    6.1, 9.7, 16.4, 14.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 0, 0.5, 1, 2, 3, 3.6, 4.1, 4.6, 5.6, 6.6, 6.6, 5.6, 3, 3.6, 2.5, 8.7, 
    11.8, 14.9, 15.9, 16.9, 15.4, 14.4, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.6, 4.1, 4.1, 3.6, 3.6, 3, 4.1, 4.1, 4.1, 2.5, 1, 1.5, 3, 3, 2, 11.8, 
    14.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2.5, 3, 3.6, 5.6, 5.6, 5.6, 5.1, 6.6, 8.7, 9.7, 12.3, 12.8, 11.8, 
    8.2, 7.7, 9.7, 9.7, 8.7, 4.1, 5.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 5.6, 7.2, 6.6, 5.6, 9.7, 10.8, 13.3, 11.8, 13.8, 15.4, 19, 21.1, 26.2, 
    26.7, 29.8, 28.3, 33.9, 39.6, 43.7, 45.8, 29.3, 17.5, 15.9, 15.9, 11.3, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.1, 7.2, 8.2, 9.2, 11.3, 10.2, 12.8, 13.3, 15.4, 19, 22.6, 27.2, 28.8, 38, 
    40.6, 40.1, 39.6, 31.4, 7.2, 9.2, 8.7, 12.3, 14.9, 11.3, 7.2, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7.7, 6.6, 9.7, 12.3, 12.8, 13.3, 14.4, 15.4, 15.4, 17.5, 20, 21.6, 22.1, 
    23.6, 29.8, 29.8, 30.8, 36.5, 40.1, 33.9, 26.7, 20.5, 18.5, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.1, 5.6, 7.2, 8.7, 12.3, 15.9, 17.5, 17.5, 20.5, 26.2, 28.3, 28.8, 28.8, 
    32.4, 36, 41.1, 36.5, 32.9, 31.4, 18, 19.5, 14.9, 13.8, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 7.7, 7.7, 8.7, 9.7, 10.2, 10.2, 9.2, 8.2, 7.7, 5.6, 3, 4.1, 4.1, 5.1, 
    7.2, 10.8, 12.3, 13.3, 19, 22.6, 14.9, 11.3, 10.8, 6.6, 4.1, 5.1, 8.2, 
    7.7, 7.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 2, 4.6, 7.7, 6.6, 6.1, 6.1, 6.6, 7.7, 9.2, 9.2, 9.2, 9.7, 10.2, 13.8, 
    12.8, 9.7, 7.7, 7.2, 6.6, 5.1, 4.6, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 2.5, 3, 6.1, 9.2, 9.7, 10.8, 11.8, 13.8, 16.9, 23.1, 25.2, 22.1, 
    17.5, 16.9, 11.3, 8.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 7.7, 11.3, 11.3, 12.3, 14.4, 15.4, 16.4, 12.3, 13.3, 12.3, 11.8, 9.7, 
    11.3, 13.3, 17.5, 14.9, 12.8, 15.4, 12.8, 10.8, 9.2, 13.8, 7.2, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 5.1, 8.2, 8.2, 8.7, 10.8, 11.3, 9.2, 9.7, 14.4, 13.8, 18.5, 16.9, 22.6, 
    33.9, 44.2, 54, 31.4, 19.5, 11.8, 13.8, 14.9, 12.3, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.6, 12.8, 17.5, 20, 21.1, 19, 16.4, 13.3, 13.8, 15.4, 15.9, 15.4, 15.4, 
    17.5, 19.5, 27.2, 25.2, 24.1, 26.2, 20, 17.5, 15.4, 15.9, 12.8, 13.8, 
    12.8, 8.7, 9.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 5.6, 10.2, 13.8, 16.9, 18.5, 21.6, 24.7, 26.7, 27.7, 24.7, 26.2, 28.3, 
    23.6, 23.1, 29.3, 34.4, 35, 48.3, 51.9, 38, 39.1, 23.6, 22.1, 19.5, 13.3, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.5, 0.5, 5.1, 0.5, 12.3, 6.1, 4.6, 5.6, 7.7, 12.8, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.5, 5.6, 5.1, 2.5, 3.6, 2, 1.5, 3.6, 4.1, 5.6, 4.6, 4.1, 5.6, 5.1, 4.6, 
    6.1, 6.1, 7.7, 10.8, 10.2, 8.2, 9.2, 9.7, 11.8, 8.7, 8.2, 8.2, 9.2, 7.2, 
    5.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 7.2, 10.8, 10.8, 12.3, 15.9, 18, 14.4, 13.8, 12.3, 11.3, 11.3, 11.8, 
    10.2, 16.9, 19, 22.6, 24.1, 25.7, 36, 45.8, 47.8, 50.9, 32.4, 27.7, 25.7, 
    18, 16.4, 10.2, 8.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1, 5.1, 6.6, 6.6, 9.2, 8.2, 8.2, 9.2, 8.7, 8.7, 10.2, 11.3, 11.3, 11.8, 
    8.2, 8.2, 10.8, 14.9, 15.9, 9.7, 9.2, 4.6, 6.6, 5.1, 5.1, 4.6, 2.5, 4.6, 
    4.1, 2.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 6.1, 6.6, 7.7, 7.7, 6.1, 5.6, 5.1, 4.6, 4.1, 4.1, 4.1, 5.1, 8.7, 13.3, 
    9.2, 7.7, 4.6, 3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  2.5, 2, 3.6, 5.1, 6.6, 4.1, 4.1, 2.5, 3, 4.6, 8.7, 16.4, 17.5, 22.1, 21.6, 
    21.1, 23.1, 28.3, 31.9, 39.1, 12.3, 9.7, 11.3, 12.3, 12.8, 10.8, 9.7, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.5, 8.2, 10.2, 9.2, 9.2, 10.2, 9.2, 9.2, 10.2, 7.2, 6.1, 8.2, 10.8, 14.4, 
    13.3, 11.8, 9.7, 11.8, 18.5, 25.2, 19.5, 15.9, 15.9, 12.3, 11.3, 15.4, 
    11.8, 12.3, 13.3, 9.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 8.7, 8.7, 9.2, 10.2, 9.7, 10.2, 7.7, 6.6, 5.1, 6.6, 6.6, 4.6, 4.6, 5.1, 
    5.6, 6.1, 6.6, 6.1, 3.6, 2.5, 3, 5.6, 7.2, 7.7, 9.2, 14.4, 15.4, 17.5, 
    23.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5, 5.1, 8.2, 9.2, 7.2, 12.3, 13.8, 13.3, 11.8, 10.2, 12.8, 17.5, 23.1, 
    26.2, 30.3, 36.5, 42.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.1, 4.6, 4.1, 7.7, 9.2, 9.2, 7.2, 3.6, 3, 3, 2.5, 2, 2.5, 3, 2, 2, 4.6, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.5, 3, 7.7, 7.2, 5.6, 5.6, 6.1, 3.6, 3, 2.5, 6.6, 6.1, 4.6, 3.6, 5.1, 5.1, 
    4.1, 4.1, 5.1, 7.2, 4.6, 8.7, 5.1, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.1, 23.6, 26.7, 35, 41.1, 34.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  7.2, 10.2, 13.3, 4.6, 1.5, 2, 4.1, 8.2, 11.3, 15.4, 18.5, 19, 26.2, 29.8, 
    42.2, 42.2, 28.3, 22.6, 14.4, 14.4, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 prTrop =
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _ ;

 tpTrop =
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _ ;

 tdTrop =
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _ ;

 wdTrop =
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _ ;

 wsTrop =
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _ ;

 prMaxW =
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _ ;

 wdMaxW =
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _ ;

 wsMaxW =
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _ ;
}
